module async_fifo_33_4_0_1_test_1 ( wr_clk, wr_reset_n, wr_en, wr_data, full, 
        afull, rd_clk, rd_reset_n, rd_en, empty, aempty, rd_data, test_si5, 
        test_si4, test_si3, test_si2, test_si1, test_so5, test_so4, test_so3, 
        test_so2, test_so1, test_se );
  input [32:0] wr_data;
  output [32:0] rd_data;
  input wr_clk, wr_reset_n, wr_en, rd_clk, rd_reset_n, rd_en, test_si5,
         test_si4, test_si3, test_si2, test_si1, test_se;
  output full, afull, empty, aempty, test_so5, test_so4, test_so3, test_so2,
         test_so1;
  wire   N45, N46, mem_3__32_, mem_3__31_, mem_3__30_, mem_3__29_, mem_3__28_,
         mem_3__27_, mem_3__26_, mem_3__25_, mem_3__24_, mem_3__23_,
         mem_3__22_, mem_3__21_, mem_3__20_, mem_3__19_, mem_3__18_,
         mem_3__17_, mem_3__16_, mem_3__15_, mem_3__14_, mem_3__13_,
         mem_3__12_, mem_3__11_, mem_3__10_, mem_3__8_, mem_3__7_, mem_3__6_,
         mem_3__5_, mem_3__4_, mem_3__3_, mem_3__2_, mem_3__1_, mem_3__0_,
         mem_2__32_, mem_2__31_, mem_2__30_, mem_2__29_, mem_2__28_,
         mem_2__27_, mem_2__26_, mem_2__25_, mem_2__24_, mem_2__23_,
         mem_2__22_, mem_2__21_, mem_2__20_, mem_2__19_, mem_2__18_,
         mem_2__17_, mem_2__16_, mem_2__15_, mem_2__14_, mem_2__13_,
         mem_2__12_, mem_2__11_, mem_2__10_, mem_2__9_, mem_2__8_, mem_2__7_,
         mem_2__6_, mem_2__5_, mem_2__4_, mem_2__3_, mem_2__2_, mem_2__1_,
         mem_2__0_, mem_1__32_, mem_1__31_, mem_1__30_, mem_1__29_, mem_1__28_,
         mem_1__26_, mem_1__25_, mem_1__24_, mem_1__23_, mem_1__22_,
         mem_1__21_, mem_1__20_, mem_1__19_, mem_1__18_, mem_1__17_,
         mem_1__16_, mem_1__15_, mem_1__14_, mem_1__13_, mem_1__12_,
         mem_1__11_, mem_1__10_, mem_1__9_, mem_1__8_, mem_1__7_, mem_1__6_,
         mem_1__5_, mem_1__4_, mem_1__3_, mem_1__2_, mem_1__1_, mem_1__0_,
         mem_0__32_, mem_0__31_, mem_0__30_, mem_0__29_, mem_0__28_,
         mem_0__27_, mem_0__26_, mem_0__25_, mem_0__24_, mem_0__23_,
         mem_0__22_, mem_0__21_, mem_0__20_, mem_0__19_, mem_0__18_,
         mem_0__17_, mem_0__16_, mem_0__15_, mem_0__14_, mem_0__13_,
         mem_0__11_, mem_0__10_, mem_0__9_, mem_0__8_, mem_0__7_, mem_0__6_,
         mem_0__5_, mem_0__4_, mem_0__3_, mem_0__2_, mem_0__1_, mem_0__0_,
         sync_wr_ptr_1_0_, n196, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n188, n189, n190, n191, n192, n193,
         n194, n195, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n614,
         n615, n616, n617, n619, n620;
  wire   [1:0] wr_ptr;
  wire   [2:0] grey_wr_ptr;
  wire   [2:0] grey_rd_ptr_dly;
  wire   [2:0] sync_rd_ptr_1;
  wire   [2:0] sync_rd_ptr_0;
  wire   [2:0] sync_wr_ptr_0;

  FD2S full_q_reg ( .D(n278), .TI(test_si2), .TE(test_se), .CP(n6), .CD(
        wr_reset_n), .Q(full), .QN(n477) );
  FD2S sync_wr_ptr_1_reg_1_ ( .D(sync_wr_ptr_0[1]), .TI(sync_wr_ptr_1_0_), 
        .TE(test_se), .CP(n26), .CD(rd_reset_n), .Q(n619), .QN(n616) );
  FD1S mem_reg_3__32_ ( .D(n314), .TI(mem_3__31_), .TE(test_se), .CP(n8), .Q(
        mem_3__32_), .QN(n510) );
  FD1S mem_reg_3__31_ ( .D(n313), .TI(mem_3__30_), .TE(test_se), .CP(n8), .Q(
        mem_3__31_), .QN(n509) );
  FD1S mem_reg_3__30_ ( .D(n312), .TI(mem_3__29_), .TE(test_se), .CP(n8), .Q(
        mem_3__30_), .QN(n508) );
  FD1S mem_reg_3__29_ ( .D(n311), .TI(mem_3__28_), .TE(test_se), .CP(n8), .Q(
        mem_3__29_), .QN(n507) );
  FD1S mem_reg_3__28_ ( .D(n310), .TI(mem_3__27_), .TE(test_se), .CP(n8), .Q(
        mem_3__28_), .QN(n506) );
  FD1S mem_reg_3__27_ ( .D(n309), .TI(mem_3__26_), .TE(test_se), .CP(n8), .Q(
        mem_3__27_), .QN(n505) );
  FD1S mem_reg_3__26_ ( .D(n308), .TI(mem_3__25_), .TE(test_se), .CP(n8), .Q(
        mem_3__26_), .QN(n504) );
  FD1S mem_reg_3__25_ ( .D(n307), .TI(mem_3__24_), .TE(test_se), .CP(n8), .Q(
        mem_3__25_), .QN(n503) );
  FD1S mem_reg_3__24_ ( .D(n306), .TI(mem_3__23_), .TE(test_se), .CP(n8), .Q(
        mem_3__24_), .QN(n502) );
  FD1S mem_reg_3__23_ ( .D(n305), .TI(mem_3__22_), .TE(test_se), .CP(n7), .Q(
        mem_3__23_), .QN(n501) );
  FD1S mem_reg_3__22_ ( .D(n304), .TI(mem_3__21_), .TE(test_se), .CP(n7), .Q(
        mem_3__22_), .QN(n500) );
  FD1S mem_reg_3__21_ ( .D(n303), .TI(mem_3__20_), .TE(test_se), .CP(n7), .Q(
        mem_3__21_), .QN(n499) );
  FD1S mem_reg_3__20_ ( .D(n302), .TI(mem_3__19_), .TE(test_se), .CP(n7), .Q(
        mem_3__20_), .QN(n498) );
  FD1S mem_reg_3__19_ ( .D(n301), .TI(mem_3__18_), .TE(test_se), .CP(n7), .Q(
        mem_3__19_), .QN(n497) );
  FD1S mem_reg_3__18_ ( .D(n300), .TI(mem_3__17_), .TE(test_se), .CP(n7), .Q(
        mem_3__18_), .QN(n496) );
  FD1S mem_reg_3__17_ ( .D(n299), .TI(mem_3__16_), .TE(test_se), .CP(n7), .Q(
        mem_3__17_), .QN(n495) );
  FD1S mem_reg_3__16_ ( .D(n298), .TI(mem_3__15_), .TE(test_se), .CP(n7), .Q(
        mem_3__16_), .QN(n494) );
  FD1S mem_reg_3__15_ ( .D(n297), .TI(mem_3__14_), .TE(test_se), .CP(n7), .Q(
        mem_3__15_), .QN(n493) );
  FD1S mem_reg_3__14_ ( .D(n296), .TI(mem_3__13_), .TE(test_se), .CP(n7), .Q(
        mem_3__14_), .QN(n492) );
  FD1S mem_reg_3__13_ ( .D(n295), .TI(mem_3__12_), .TE(test_se), .CP(n7), .Q(
        mem_3__13_), .QN(n491) );
  FD1S mem_reg_3__12_ ( .D(n294), .TI(mem_3__11_), .TE(test_se), .CP(n7), .Q(
        mem_3__12_), .QN(n490) );
  FD1S mem_reg_3__11_ ( .D(n293), .TI(mem_3__10_), .TE(test_se), .CP(n6), .Q(
        mem_3__11_), .QN(n489) );
  FD1S mem_reg_3__10_ ( .D(n292), .TI(test_si5), .TE(test_se), .CP(n6), .Q(
        mem_3__10_), .QN(n488) );
  FD1S mem_reg_3__9_ ( .D(n291), .TI(mem_3__8_), .TE(test_se), .CP(n6), .Q(
        test_so4), .QN(n487) );
  FD1S mem_reg_3__8_ ( .D(n290), .TI(mem_3__7_), .TE(test_se), .CP(n6), .Q(
        mem_3__8_), .QN(n486) );
  FD1S mem_reg_3__7_ ( .D(n289), .TI(mem_3__6_), .TE(test_se), .CP(n6), .Q(
        mem_3__7_), .QN(n485) );
  FD1S mem_reg_3__6_ ( .D(n288), .TI(mem_3__5_), .TE(test_se), .CP(n6), .Q(
        mem_3__6_), .QN(n484) );
  FD1S mem_reg_3__5_ ( .D(n287), .TI(mem_3__4_), .TE(test_se), .CP(n6), .Q(
        mem_3__5_), .QN(n483) );
  FD1S mem_reg_3__4_ ( .D(n286), .TI(mem_3__3_), .TE(test_se), .CP(n6), .Q(
        mem_3__4_), .QN(n482) );
  FD1S mem_reg_3__3_ ( .D(n285), .TI(mem_3__2_), .TE(test_se), .CP(n6), .Q(
        mem_3__3_), .QN(n481) );
  FD1S mem_reg_3__2_ ( .D(n284), .TI(mem_3__1_), .TE(test_se), .CP(n6), .Q(
        mem_3__2_), .QN(n480) );
  FD1S mem_reg_3__1_ ( .D(n283), .TI(mem_3__0_), .TE(test_se), .CP(n6), .Q(
        mem_3__1_), .QN(n479) );
  FD1S mem_reg_3__0_ ( .D(n315), .TI(mem_2__32_), .TE(test_se), .CP(n8), .Q(
        mem_3__0_), .QN(n511) );
  FD1S mem_reg_2__32_ ( .D(n347), .TI(mem_2__31_), .TE(test_se), .CP(n11), .Q(
        mem_2__32_), .QN(n543) );
  FD1S mem_reg_2__31_ ( .D(n346), .TI(mem_2__30_), .TE(test_se), .CP(n11), .Q(
        mem_2__31_), .QN(n542) );
  FD1S mem_reg_2__30_ ( .D(n345), .TI(mem_2__29_), .TE(test_se), .CP(n11), .Q(
        mem_2__30_), .QN(n541) );
  FD1S mem_reg_2__29_ ( .D(n344), .TI(mem_2__28_), .TE(test_se), .CP(n11), .Q(
        mem_2__29_), .QN(n540) );
  FD1S mem_reg_2__28_ ( .D(n343), .TI(mem_2__27_), .TE(test_se), .CP(n11), .Q(
        mem_2__28_), .QN(n539) );
  FD1S mem_reg_2__27_ ( .D(n342), .TI(mem_2__26_), .TE(test_se), .CP(n11), .Q(
        mem_2__27_), .QN(n538) );
  FD1S mem_reg_2__26_ ( .D(n341), .TI(mem_2__25_), .TE(test_se), .CP(n10), .Q(
        mem_2__26_), .QN(n537) );
  FD1S mem_reg_2__25_ ( .D(n340), .TI(mem_2__24_), .TE(test_se), .CP(n10), .Q(
        mem_2__25_), .QN(n536) );
  FD1S mem_reg_2__24_ ( .D(n339), .TI(mem_2__23_), .TE(test_se), .CP(n10), .Q(
        mem_2__24_), .QN(n535) );
  FD1S mem_reg_2__23_ ( .D(n338), .TI(mem_2__22_), .TE(test_se), .CP(n10), .Q(
        mem_2__23_), .QN(n534) );
  FD1S mem_reg_2__22_ ( .D(n337), .TI(mem_2__21_), .TE(test_se), .CP(n10), .Q(
        mem_2__22_), .QN(n533) );
  FD1S mem_reg_2__21_ ( .D(n336), .TI(mem_2__20_), .TE(test_se), .CP(n10), .Q(
        mem_2__21_), .QN(n532) );
  FD1S mem_reg_2__20_ ( .D(n335), .TI(mem_2__19_), .TE(test_se), .CP(n10), .Q(
        mem_2__20_), .QN(n531) );
  FD1S mem_reg_2__19_ ( .D(n334), .TI(mem_2__18_), .TE(test_se), .CP(n10), .Q(
        mem_2__19_), .QN(n530) );
  FD1S mem_reg_2__18_ ( .D(n333), .TI(mem_2__17_), .TE(test_se), .CP(n10), .Q(
        mem_2__18_), .QN(n529) );
  FD1S mem_reg_2__17_ ( .D(n332), .TI(mem_2__16_), .TE(test_se), .CP(n10), .Q(
        mem_2__17_), .QN(n528) );
  FD1S mem_reg_2__16_ ( .D(n331), .TI(mem_2__15_), .TE(test_se), .CP(n10), .Q(
        mem_2__16_), .QN(n527) );
  FD1S mem_reg_2__15_ ( .D(n330), .TI(mem_2__14_), .TE(test_se), .CP(n10), .Q(
        mem_2__15_), .QN(n526) );
  FD1S mem_reg_2__14_ ( .D(n329), .TI(mem_2__13_), .TE(test_se), .CP(n9), .Q(
        mem_2__14_), .QN(n525) );
  FD1S mem_reg_2__13_ ( .D(n328), .TI(mem_2__12_), .TE(test_se), .CP(n9), .Q(
        mem_2__13_), .QN(n524) );
  FD1S mem_reg_2__12_ ( .D(n327), .TI(mem_2__11_), .TE(test_se), .CP(n9), .Q(
        mem_2__12_), .QN(n523) );
  FD1S mem_reg_2__11_ ( .D(n326), .TI(mem_2__10_), .TE(test_se), .CP(n9), .Q(
        mem_2__11_), .QN(n522) );
  FD1S mem_reg_2__10_ ( .D(n325), .TI(mem_2__9_), .TE(test_se), .CP(n9), .Q(
        mem_2__10_), .QN(n521) );
  FD1S mem_reg_2__9_ ( .D(n324), .TI(mem_2__8_), .TE(test_se), .CP(n9), .Q(
        mem_2__9_), .QN(n520) );
  FD1S mem_reg_2__8_ ( .D(n323), .TI(mem_2__7_), .TE(test_se), .CP(n9), .Q(
        mem_2__8_), .QN(n519) );
  FD1S mem_reg_2__7_ ( .D(n322), .TI(mem_2__6_), .TE(test_se), .CP(n9), .Q(
        mem_2__7_), .QN(n518) );
  FD1S mem_reg_2__6_ ( .D(n321), .TI(mem_2__5_), .TE(test_se), .CP(n9), .Q(
        mem_2__6_), .QN(n517) );
  FD1S mem_reg_2__5_ ( .D(n320), .TI(mem_2__4_), .TE(test_se), .CP(n9), .Q(
        mem_2__5_), .QN(n516) );
  FD1S mem_reg_2__4_ ( .D(n319), .TI(mem_2__3_), .TE(test_se), .CP(n9), .Q(
        mem_2__4_), .QN(n515) );
  FD1S mem_reg_2__3_ ( .D(n318), .TI(mem_2__2_), .TE(test_se), .CP(n9), .Q(
        mem_2__3_), .QN(n514) );
  FD1S mem_reg_2__2_ ( .D(n317), .TI(mem_2__1_), .TE(test_se), .CP(n8), .Q(
        mem_2__2_), .QN(n513) );
  FD1S mem_reg_2__1_ ( .D(n316), .TI(mem_2__0_), .TE(test_se), .CP(n8), .Q(
        mem_2__1_), .QN(n512) );
  FD1S mem_reg_2__0_ ( .D(n348), .TI(mem_1__32_), .TE(test_se), .CP(n11), .Q(
        mem_2__0_), .QN(n544) );
  FD1S mem_reg_1__32_ ( .D(n380), .TI(mem_1__31_), .TE(test_se), .CP(n14), .Q(
        mem_1__32_), .QN(n576) );
  FD1S mem_reg_1__31_ ( .D(n379), .TI(mem_1__30_), .TE(test_se), .CP(n14), .Q(
        mem_1__31_), .QN(n575) );
  FD1S mem_reg_1__30_ ( .D(n378), .TI(mem_1__29_), .TE(test_se), .CP(n14), .Q(
        mem_1__30_), .QN(n574) );
  FD1S mem_reg_1__29_ ( .D(n377), .TI(mem_1__28_), .TE(test_se), .CP(n13), .Q(
        mem_1__29_), .QN(n573) );
  FD1S mem_reg_1__28_ ( .D(n376), .TI(test_si4), .TE(test_se), .CP(n13), .Q(
        mem_1__28_), .QN(n572) );
  FD1S mem_reg_1__27_ ( .D(n375), .TI(mem_1__26_), .TE(test_se), .CP(n13), .Q(
        test_so3), .QN(n571) );
  FD1S mem_reg_1__26_ ( .D(n374), .TI(mem_1__25_), .TE(test_se), .CP(n13), .Q(
        mem_1__26_), .QN(n570) );
  FD1S mem_reg_1__25_ ( .D(n373), .TI(mem_1__24_), .TE(test_se), .CP(n13), .Q(
        mem_1__25_), .QN(n569) );
  FD1S mem_reg_1__24_ ( .D(n372), .TI(mem_1__23_), .TE(test_se), .CP(n13), .Q(
        mem_1__24_), .QN(n568) );
  FD1S mem_reg_1__23_ ( .D(n371), .TI(mem_1__22_), .TE(test_se), .CP(n13), .Q(
        mem_1__23_), .QN(n567) );
  FD1S mem_reg_1__22_ ( .D(n370), .TI(mem_1__21_), .TE(test_se), .CP(n13), .Q(
        mem_1__22_), .QN(n566) );
  FD1S mem_reg_1__21_ ( .D(n369), .TI(mem_1__20_), .TE(test_se), .CP(n13), .Q(
        mem_1__21_), .QN(n565) );
  FD1S mem_reg_1__20_ ( .D(n368), .TI(mem_1__19_), .TE(test_se), .CP(n13), .Q(
        mem_1__20_), .QN(n564) );
  FD1S mem_reg_1__19_ ( .D(n367), .TI(mem_1__18_), .TE(test_se), .CP(n13), .Q(
        mem_1__19_), .QN(n563) );
  FD1S mem_reg_1__18_ ( .D(n366), .TI(mem_1__17_), .TE(test_se), .CP(n13), .Q(
        mem_1__18_), .QN(n562) );
  FD1S mem_reg_1__17_ ( .D(n365), .TI(mem_1__16_), .TE(test_se), .CP(n12), .Q(
        mem_1__17_), .QN(n561) );
  FD1S mem_reg_1__16_ ( .D(n364), .TI(mem_1__15_), .TE(test_se), .CP(n12), .Q(
        mem_1__16_), .QN(n560) );
  FD1S mem_reg_1__15_ ( .D(n363), .TI(mem_1__14_), .TE(test_se), .CP(n12), .Q(
        mem_1__15_), .QN(n559) );
  FD1S mem_reg_1__14_ ( .D(n362), .TI(mem_1__13_), .TE(test_se), .CP(n12), .Q(
        mem_1__14_), .QN(n558) );
  FD1S mem_reg_1__13_ ( .D(n361), .TI(mem_1__12_), .TE(test_se), .CP(n12), .Q(
        mem_1__13_), .QN(n557) );
  FD1S mem_reg_1__12_ ( .D(n360), .TI(mem_1__11_), .TE(test_se), .CP(n12), .Q(
        mem_1__12_), .QN(n556) );
  FD1S mem_reg_1__11_ ( .D(n359), .TI(mem_1__10_), .TE(test_se), .CP(n12), .Q(
        mem_1__11_), .QN(n555) );
  FD1S mem_reg_1__10_ ( .D(n358), .TI(mem_1__9_), .TE(test_se), .CP(n12), .Q(
        mem_1__10_), .QN(n554) );
  FD1S mem_reg_1__9_ ( .D(n357), .TI(mem_1__8_), .TE(test_se), .CP(n12), .Q(
        mem_1__9_), .QN(n553) );
  FD1S mem_reg_1__8_ ( .D(n356), .TI(mem_1__7_), .TE(test_se), .CP(n12), .Q(
        mem_1__8_), .QN(n552) );
  FD1S mem_reg_1__7_ ( .D(n355), .TI(mem_1__6_), .TE(test_se), .CP(n12), .Q(
        mem_1__7_), .QN(n551) );
  FD1S mem_reg_1__6_ ( .D(n354), .TI(mem_1__5_), .TE(test_se), .CP(n12), .Q(
        mem_1__6_), .QN(n550) );
  FD1S mem_reg_1__5_ ( .D(n353), .TI(mem_1__4_), .TE(test_se), .CP(n11), .Q(
        mem_1__5_), .QN(n549) );
  FD1S mem_reg_1__4_ ( .D(n352), .TI(mem_1__3_), .TE(test_se), .CP(n11), .Q(
        mem_1__4_), .QN(n548) );
  FD1S mem_reg_1__3_ ( .D(n351), .TI(mem_1__2_), .TE(test_se), .CP(n11), .Q(
        mem_1__3_), .QN(n547) );
  FD1S mem_reg_1__2_ ( .D(n350), .TI(mem_1__1_), .TE(test_se), .CP(n11), .Q(
        mem_1__2_), .QN(n546) );
  FD1S mem_reg_1__1_ ( .D(n349), .TI(mem_1__0_), .TE(test_se), .CP(n11), .Q(
        mem_1__1_), .QN(n545) );
  FD1S mem_reg_1__0_ ( .D(n381), .TI(mem_0__32_), .TE(test_se), .CP(n14), .Q(
        mem_1__0_), .QN(n577) );
  FD1S mem_reg_0__32_ ( .D(n413), .TI(mem_0__31_), .TE(test_se), .CP(n16), .Q(
        mem_0__32_), .QN(n609) );
  FD1S mem_reg_0__31_ ( .D(n412), .TI(mem_0__30_), .TE(test_se), .CP(n16), .Q(
        mem_0__31_), .QN(n608) );
  FD1S mem_reg_0__30_ ( .D(n411), .TI(mem_0__29_), .TE(test_se), .CP(n16), .Q(
        mem_0__30_), .QN(n607) );
  FD1S mem_reg_0__29_ ( .D(n410), .TI(mem_0__28_), .TE(test_se), .CP(n16), .Q(
        mem_0__29_), .QN(n606) );
  FD1S mem_reg_0__28_ ( .D(n409), .TI(mem_0__27_), .TE(test_se), .CP(n16), .Q(
        mem_0__28_), .QN(n605) );
  FD1S mem_reg_0__27_ ( .D(n408), .TI(mem_0__26_), .TE(test_se), .CP(n16), .Q(
        mem_0__27_), .QN(n604) );
  FD1S mem_reg_0__26_ ( .D(n407), .TI(mem_0__25_), .TE(test_se), .CP(n16), .Q(
        mem_0__26_), .QN(n603) );
  FD1S mem_reg_0__25_ ( .D(n406), .TI(mem_0__24_), .TE(test_se), .CP(n16), .Q(
        mem_0__25_), .QN(n602) );
  FD1S mem_reg_0__24_ ( .D(n405), .TI(mem_0__23_), .TE(test_se), .CP(n16), .Q(
        mem_0__24_), .QN(n601) );
  FD1S mem_reg_0__23_ ( .D(n404), .TI(mem_0__22_), .TE(test_se), .CP(n16), .Q(
        mem_0__23_), .QN(n600) );
  FD1S mem_reg_0__22_ ( .D(n403), .TI(mem_0__21_), .TE(test_se), .CP(n16), .Q(
        mem_0__22_), .QN(n599) );
  FD1S mem_reg_0__21_ ( .D(n402), .TI(mem_0__20_), .TE(test_se), .CP(n16), .Q(
        mem_0__21_), .QN(n598) );
  FD1S mem_reg_0__20_ ( .D(n401), .TI(mem_0__19_), .TE(test_se), .CP(n15), .Q(
        mem_0__20_), .QN(n597) );
  FD1S mem_reg_0__19_ ( .D(n400), .TI(mem_0__18_), .TE(test_se), .CP(n15), .Q(
        mem_0__19_), .QN(n596) );
  FD1S mem_reg_0__18_ ( .D(n399), .TI(mem_0__17_), .TE(test_se), .CP(n15), .Q(
        mem_0__18_), .QN(n595) );
  FD1S mem_reg_0__17_ ( .D(n398), .TI(mem_0__16_), .TE(test_se), .CP(n15), .Q(
        mem_0__17_), .QN(n594) );
  FD1S mem_reg_0__16_ ( .D(n397), .TI(mem_0__15_), .TE(test_se), .CP(n15), .Q(
        mem_0__16_), .QN(n593) );
  FD1S mem_reg_0__15_ ( .D(n396), .TI(mem_0__14_), .TE(test_se), .CP(n15), .Q(
        mem_0__15_), .QN(n592) );
  FD1S mem_reg_0__14_ ( .D(n395), .TI(mem_0__13_), .TE(test_se), .CP(n15), .Q(
        mem_0__14_), .QN(n591) );
  FD1S mem_reg_0__13_ ( .D(n394), .TI(test_si3), .TE(test_se), .CP(n15), .Q(
        mem_0__13_), .QN(n590) );
  FD1S mem_reg_0__12_ ( .D(n393), .TI(mem_0__11_), .TE(test_se), .CP(n15), .Q(
        test_so2), .QN(n589) );
  FD1S mem_reg_0__11_ ( .D(n392), .TI(mem_0__10_), .TE(test_se), .CP(n15), .Q(
        mem_0__11_), .QN(n588) );
  FD1S mem_reg_0__10_ ( .D(n391), .TI(mem_0__9_), .TE(test_se), .CP(n15), .Q(
        mem_0__10_), .QN(n587) );
  FD1S mem_reg_0__9_ ( .D(n390), .TI(mem_0__8_), .TE(test_se), .CP(n15), .Q(
        mem_0__9_), .QN(n586) );
  FD1S mem_reg_0__8_ ( .D(n389), .TI(mem_0__7_), .TE(test_se), .CP(n14), .Q(
        mem_0__8_), .QN(n585) );
  FD1S mem_reg_0__7_ ( .D(n388), .TI(mem_0__6_), .TE(test_se), .CP(n14), .Q(
        mem_0__7_), .QN(n584) );
  FD1S mem_reg_0__6_ ( .D(n387), .TI(mem_0__5_), .TE(test_se), .CP(n14), .Q(
        mem_0__6_), .QN(n583) );
  FD1S mem_reg_0__5_ ( .D(n386), .TI(mem_0__4_), .TE(test_se), .CP(n14), .Q(
        mem_0__5_), .QN(n582) );
  FD1S mem_reg_0__4_ ( .D(n385), .TI(mem_0__3_), .TE(test_se), .CP(n14), .Q(
        mem_0__4_), .QN(n581) );
  FD1S mem_reg_0__3_ ( .D(n384), .TI(mem_0__2_), .TE(test_se), .CP(n14), .Q(
        mem_0__3_), .QN(n580) );
  FD1S mem_reg_0__2_ ( .D(n383), .TI(mem_0__1_), .TE(test_se), .CP(n14), .Q(
        mem_0__2_), .QN(n579) );
  FD1S mem_reg_0__1_ ( .D(n382), .TI(mem_0__0_), .TE(test_se), .CP(n14), .Q(
        mem_0__1_), .QN(n578) );
  FD1S mem_reg_0__0_ ( .D(n414), .TI(grey_wr_ptr[2]), .TE(test_se), .CP(n17), 
        .Q(mem_0__0_), .QN(n610) );
  FD2S grey_wr_ptr_reg_2_ ( .D(n281), .TI(grey_wr_ptr[1]), .TE(test_se), .CP(
        n5), .CD(wr_reset_n), .Q(grey_wr_ptr[2]), .QN(n478) );
  FD2S grey_rd_ptr_reg_1_ ( .D(n416), .TI(grey_rd_ptr_dly[0]), .TE(test_se), 
        .CP(n26), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[1]), .QN(n611) );
  FD2S grey_rd_ptr_reg_2_ ( .D(n418), .TI(grey_rd_ptr_dly[1]), .TE(test_se), 
        .CP(n26), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[2]), .QN(n612) );
  FD2S rd_ptr_reg_2_ ( .D(n419), .TI(N46), .TE(test_se), .CP(n26), .CD(
        rd_reset_n), .Q(n620), .QN(n3) );
  FD2S grey_wr_ptr_reg_1_ ( .D(n279), .TI(grey_wr_ptr[0]), .TE(test_se), .CP(
        n5), .CD(wr_reset_n), .Q(grey_wr_ptr[1]) );
  FD2S sync_rd_ptr_1_reg_0_ ( .D(sync_rd_ptr_0[0]), .TI(sync_rd_ptr_0[2]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[0]) );
  FD2S sync_rd_ptr_1_reg_1_ ( .D(sync_rd_ptr_0[1]), .TI(sync_rd_ptr_1[0]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[1]), .QN(n614) );
  FD2S sync_wr_ptr_1_reg_0_ ( .D(sync_wr_ptr_0[0]), .TI(sync_wr_ptr_0[2]), 
        .TE(test_se), .CP(n26), .CD(rd_reset_n), .Q(sync_wr_ptr_1_0_) );
  FD2S wr_ptr_reg_2_ ( .D(n282), .TI(wr_ptr[1]), .TE(test_se), .CP(n5), .CD(
        wr_reset_n), .Q(test_so5), .QN(n2) );
  FD2S grey_wr_ptr_reg_0_ ( .D(n280), .TI(full), .TE(test_se), .CP(n5), .CD(
        wr_reset_n), .Q(grey_wr_ptr[0]) );
  FD2S grey_rd_ptr_reg_0_ ( .D(n417), .TI(test_si1), .TE(test_se), .CP(n26), 
        .CD(rd_reset_n), .Q(grey_rd_ptr_dly[0]) );
  FD2S sync_rd_ptr_1_reg_2_ ( .D(sync_rd_ptr_0[2]), .TI(sync_rd_ptr_1[1]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[2]) );
  FD2S sync_wr_ptr_1_reg_2_ ( .D(sync_wr_ptr_0[2]), .TI(n619), .TE(test_se), 
        .CP(n26), .CD(rd_reset_n), .Q(test_so1) );
  FD2S wr_ptr_reg_1_ ( .D(n415), .TI(wr_ptr[0]), .TE(test_se), .CP(n5), .CD(
        wr_reset_n), .Q(wr_ptr[1]), .QN(n1) );
  FD2S rd_ptr_reg_0_ ( .D(n421), .TI(grey_rd_ptr_dly[2]), .TE(test_se), .CP(
        n26), .CD(rd_reset_n), .Q(N45), .QN(n615) );
  FD2S rd_ptr_reg_1_ ( .D(n420), .TI(N45), .TE(test_se), .CP(n26), .CD(
        rd_reset_n), .Q(N46), .QN(n196) );
  FD2S wr_ptr_reg_0_ ( .D(n617), .TI(sync_rd_ptr_1[2]), .TE(test_se), .CP(n5), 
        .CD(wr_reset_n), .Q(wr_ptr[0]), .QN(n4) );
  FD2S sync_wr_ptr_0_reg_2_ ( .D(grey_wr_ptr[2]), .TI(sync_wr_ptr_0[1]), .TE(
        test_se), .CP(n26), .CD(rd_reset_n), .Q(sync_wr_ptr_0[2]) );
  FD2S sync_wr_ptr_0_reg_1_ ( .D(grey_wr_ptr[1]), .TI(sync_wr_ptr_0[0]), .TE(
        test_se), .CP(n26), .CD(rd_reset_n), .Q(sync_wr_ptr_0[1]) );
  FD2S sync_wr_ptr_0_reg_0_ ( .D(grey_wr_ptr[0]), .TI(n620), .TE(test_se), 
        .CP(n26), .CD(rd_reset_n), .Q(sync_wr_ptr_0[0]) );
  FD2S sync_rd_ptr_0_reg_0_ ( .D(grey_rd_ptr_dly[0]), .TI(mem_3__32_), .TE(
        test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[0]) );
  FD2S sync_rd_ptr_0_reg_1_ ( .D(grey_rd_ptr_dly[1]), .TI(sync_rd_ptr_0[0]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[1]) );
  FD2S sync_rd_ptr_0_reg_2_ ( .D(grey_rd_ptr_dly[2]), .TI(sync_rd_ptr_0[1]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[2]) );
  IVP U160 ( .A(n18), .Z(n15) );
  IVP U161 ( .A(n18), .Z(n16) );
  IVP U162 ( .A(n19), .Z(n12) );
  IVP U163 ( .A(n19), .Z(n13) );
  IVP U164 ( .A(n19), .Z(n14) );
  IVP U165 ( .A(n20), .Z(n9) );
  IVP U166 ( .A(n20), .Z(n10) );
  IVP U167 ( .A(n20), .Z(n11) );
  IVP U168 ( .A(n21), .Z(n6) );
  IVP U169 ( .A(n21), .Z(n7) );
  IVP U170 ( .A(n21), .Z(n8) );
  IVP U171 ( .A(n18), .Z(n17) );
  IVP U172 ( .A(n24), .Z(n18) );
  IVP U173 ( .A(n24), .Z(n19) );
  IVP U174 ( .A(n23), .Z(n20) );
  IVP U175 ( .A(n23), .Z(n21) );
  IVP U176 ( .A(n22), .Z(n5) );
  IVP U177 ( .A(n23), .Z(n22) );
  IVP U178 ( .A(n25), .Z(n23) );
  IVP U179 ( .A(n25), .Z(n24) );
  IVP U180 ( .A(wr_clk), .Z(n25) );
  IVP U181 ( .A(n27), .Z(n26) );
  IVP U182 ( .A(rd_clk), .Z(n27) );
  NR2 U183 ( .A(n196), .B(N45), .Z(n251) );
  NR2 U184 ( .A(n196), .B(n615), .Z(n250) );
  AO2 U185 ( .A(mem_2__0_), .B(n251), .C(mem_3__0_), .D(n250), .Z(n29) );
  NR2 U186 ( .A(N45), .B(N46), .Z(n253) );
  NR2 U187 ( .A(n615), .B(N46), .Z(n252) );
  AO2 U188 ( .A(mem_0__0_), .B(n253), .C(mem_1__0_), .D(n252), .Z(n28) );
  ND2 U189 ( .A(n29), .B(n28), .Z(rd_data[0]) );
  AO2 U190 ( .A(mem_2__1_), .B(n251), .C(mem_3__1_), .D(n250), .Z(n188) );
  AO2 U191 ( .A(mem_0__1_), .B(n253), .C(mem_1__1_), .D(n252), .Z(n30) );
  ND2 U192 ( .A(n188), .B(n30), .Z(rd_data[1]) );
  AO2 U193 ( .A(mem_2__2_), .B(n251), .C(mem_3__2_), .D(n250), .Z(n190) );
  AO2 U194 ( .A(mem_0__2_), .B(n253), .C(mem_1__2_), .D(n252), .Z(n189) );
  ND2 U195 ( .A(n190), .B(n189), .Z(rd_data[2]) );
  AO2 U196 ( .A(mem_2__3_), .B(n251), .C(mem_3__3_), .D(n250), .Z(n192) );
  AO2 U197 ( .A(mem_0__3_), .B(n253), .C(mem_1__3_), .D(n252), .Z(n191) );
  ND2 U198 ( .A(n192), .B(n191), .Z(rd_data[3]) );
  AO2 U199 ( .A(mem_2__4_), .B(n251), .C(mem_3__4_), .D(n250), .Z(n194) );
  AO2 U200 ( .A(mem_0__4_), .B(n253), .C(mem_1__4_), .D(n252), .Z(n193) );
  ND2 U201 ( .A(n194), .B(n193), .Z(rd_data[4]) );
  AO2 U202 ( .A(mem_2__5_), .B(n251), .C(mem_3__5_), .D(n250), .Z(n197) );
  AO2 U203 ( .A(mem_0__5_), .B(n253), .C(mem_1__5_), .D(n252), .Z(n195) );
  ND2 U204 ( .A(n197), .B(n195), .Z(rd_data[5]) );
  AO2 U205 ( .A(mem_2__6_), .B(n251), .C(mem_3__6_), .D(n250), .Z(n199) );
  AO2 U206 ( .A(mem_0__6_), .B(n253), .C(mem_1__6_), .D(n252), .Z(n198) );
  ND2 U207 ( .A(n199), .B(n198), .Z(rd_data[6]) );
  AO2 U208 ( .A(mem_2__7_), .B(n251), .C(mem_3__7_), .D(n250), .Z(n201) );
  AO2 U209 ( .A(mem_0__7_), .B(n253), .C(mem_1__7_), .D(n252), .Z(n200) );
  ND2 U210 ( .A(n201), .B(n200), .Z(rd_data[7]) );
  AO2 U211 ( .A(mem_2__8_), .B(n251), .C(mem_3__8_), .D(n250), .Z(n203) );
  AO2 U212 ( .A(mem_0__8_), .B(n253), .C(mem_1__8_), .D(n252), .Z(n202) );
  ND2 U213 ( .A(n203), .B(n202), .Z(rd_data[8]) );
  AO2 U214 ( .A(mem_2__9_), .B(n251), .C(test_so4), .D(n250), .Z(n205) );
  AO2 U215 ( .A(mem_0__9_), .B(n253), .C(mem_1__9_), .D(n252), .Z(n204) );
  ND2 U216 ( .A(n205), .B(n204), .Z(rd_data[9]) );
  AO2 U217 ( .A(mem_2__10_), .B(n251), .C(mem_3__10_), .D(n250), .Z(n207) );
  AO2 U218 ( .A(mem_0__10_), .B(n253), .C(mem_1__10_), .D(n252), .Z(n206) );
  ND2 U219 ( .A(n207), .B(n206), .Z(rd_data[10]) );
  AO2 U220 ( .A(mem_2__11_), .B(n251), .C(mem_3__11_), .D(n250), .Z(n209) );
  AO2 U221 ( .A(mem_0__11_), .B(n253), .C(mem_1__11_), .D(n252), .Z(n208) );
  ND2 U222 ( .A(n209), .B(n208), .Z(rd_data[11]) );
  AO2 U223 ( .A(mem_2__12_), .B(n251), .C(mem_3__12_), .D(n250), .Z(n211) );
  AO2 U224 ( .A(test_so2), .B(n253), .C(mem_1__12_), .D(n252), .Z(n210) );
  ND2 U225 ( .A(n211), .B(n210), .Z(rd_data[12]) );
  AO2 U226 ( .A(mem_2__13_), .B(n251), .C(mem_3__13_), .D(n250), .Z(n213) );
  AO2 U227 ( .A(mem_0__13_), .B(n253), .C(mem_1__13_), .D(n252), .Z(n212) );
  ND2 U228 ( .A(n213), .B(n212), .Z(rd_data[13]) );
  AO2 U229 ( .A(mem_2__14_), .B(n251), .C(mem_3__14_), .D(n250), .Z(n215) );
  AO2 U230 ( .A(mem_0__14_), .B(n253), .C(mem_1__14_), .D(n252), .Z(n214) );
  ND2 U231 ( .A(n215), .B(n214), .Z(rd_data[14]) );
  AO2 U232 ( .A(mem_2__15_), .B(n251), .C(mem_3__15_), .D(n250), .Z(n217) );
  AO2 U233 ( .A(mem_0__15_), .B(n253), .C(mem_1__15_), .D(n252), .Z(n216) );
  ND2 U234 ( .A(n217), .B(n216), .Z(rd_data[15]) );
  AO2 U235 ( .A(mem_2__16_), .B(n251), .C(mem_3__16_), .D(n250), .Z(n219) );
  AO2 U236 ( .A(mem_0__16_), .B(n253), .C(mem_1__16_), .D(n252), .Z(n218) );
  ND2 U237 ( .A(n219), .B(n218), .Z(rd_data[16]) );
  AO2 U238 ( .A(mem_2__17_), .B(n251), .C(mem_3__17_), .D(n250), .Z(n221) );
  AO2 U239 ( .A(mem_0__17_), .B(n253), .C(mem_1__17_), .D(n252), .Z(n220) );
  ND2 U240 ( .A(n221), .B(n220), .Z(rd_data[17]) );
  AO2 U241 ( .A(mem_2__18_), .B(n251), .C(mem_3__18_), .D(n250), .Z(n223) );
  AO2 U242 ( .A(mem_0__18_), .B(n253), .C(mem_1__18_), .D(n252), .Z(n222) );
  ND2 U243 ( .A(n223), .B(n222), .Z(rd_data[18]) );
  AO2 U244 ( .A(mem_2__19_), .B(n251), .C(mem_3__19_), .D(n250), .Z(n225) );
  AO2 U245 ( .A(mem_0__19_), .B(n253), .C(mem_1__19_), .D(n252), .Z(n224) );
  ND2 U246 ( .A(n225), .B(n224), .Z(rd_data[19]) );
  AO2 U247 ( .A(mem_2__20_), .B(n251), .C(mem_3__20_), .D(n250), .Z(n227) );
  AO2 U248 ( .A(mem_0__20_), .B(n253), .C(mem_1__20_), .D(n252), .Z(n226) );
  ND2 U249 ( .A(n227), .B(n226), .Z(rd_data[20]) );
  AO2 U250 ( .A(mem_2__21_), .B(n251), .C(mem_3__21_), .D(n250), .Z(n229) );
  AO2 U251 ( .A(mem_0__21_), .B(n253), .C(mem_1__21_), .D(n252), .Z(n228) );
  ND2 U252 ( .A(n229), .B(n228), .Z(rd_data[21]) );
  AO2 U253 ( .A(mem_2__22_), .B(n251), .C(mem_3__22_), .D(n250), .Z(n231) );
  AO2 U254 ( .A(mem_0__22_), .B(n253), .C(mem_1__22_), .D(n252), .Z(n230) );
  ND2 U255 ( .A(n231), .B(n230), .Z(rd_data[22]) );
  AO2 U256 ( .A(mem_2__23_), .B(n251), .C(mem_3__23_), .D(n250), .Z(n233) );
  AO2 U257 ( .A(mem_0__23_), .B(n253), .C(mem_1__23_), .D(n252), .Z(n232) );
  ND2 U258 ( .A(n233), .B(n232), .Z(rd_data[23]) );
  AO2 U259 ( .A(mem_2__24_), .B(n251), .C(mem_3__24_), .D(n250), .Z(n235) );
  AO2 U260 ( .A(mem_0__24_), .B(n253), .C(mem_1__24_), .D(n252), .Z(n234) );
  ND2 U261 ( .A(n235), .B(n234), .Z(rd_data[24]) );
  AO2 U262 ( .A(mem_2__25_), .B(n251), .C(mem_3__25_), .D(n250), .Z(n237) );
  AO2 U263 ( .A(mem_0__25_), .B(n253), .C(mem_1__25_), .D(n252), .Z(n236) );
  ND2 U264 ( .A(n237), .B(n236), .Z(rd_data[25]) );
  AO2 U265 ( .A(mem_2__26_), .B(n251), .C(mem_3__26_), .D(n250), .Z(n239) );
  AO2 U266 ( .A(mem_0__26_), .B(n253), .C(mem_1__26_), .D(n252), .Z(n238) );
  ND2 U267 ( .A(n239), .B(n238), .Z(rd_data[26]) );
  AO2 U268 ( .A(mem_2__27_), .B(n251), .C(mem_3__27_), .D(n250), .Z(n241) );
  AO2 U269 ( .A(mem_0__27_), .B(n253), .C(test_so3), .D(n252), .Z(n240) );
  ND2 U270 ( .A(n241), .B(n240), .Z(rd_data[27]) );
  AO2 U271 ( .A(mem_2__28_), .B(n251), .C(mem_3__28_), .D(n250), .Z(n243) );
  AO2 U272 ( .A(mem_0__28_), .B(n253), .C(mem_1__28_), .D(n252), .Z(n242) );
  ND2 U273 ( .A(n243), .B(n242), .Z(rd_data[28]) );
  AO2 U274 ( .A(mem_2__29_), .B(n251), .C(mem_3__29_), .D(n250), .Z(n245) );
  AO2 U275 ( .A(mem_0__29_), .B(n253), .C(mem_1__29_), .D(n252), .Z(n244) );
  ND2 U276 ( .A(n245), .B(n244), .Z(rd_data[29]) );
  AO2 U277 ( .A(mem_2__30_), .B(n251), .C(mem_3__30_), .D(n250), .Z(n247) );
  AO2 U278 ( .A(mem_0__30_), .B(n253), .C(mem_1__30_), .D(n252), .Z(n246) );
  ND2 U279 ( .A(n247), .B(n246), .Z(rd_data[30]) );
  AO2 U280 ( .A(mem_2__31_), .B(n251), .C(mem_3__31_), .D(n250), .Z(n249) );
  AO2 U281 ( .A(mem_0__31_), .B(n253), .C(mem_1__31_), .D(n252), .Z(n248) );
  ND2 U282 ( .A(n249), .B(n248), .Z(rd_data[31]) );
  AO2 U283 ( .A(mem_2__32_), .B(n251), .C(mem_3__32_), .D(n250), .Z(n255) );
  AO2 U284 ( .A(mem_0__32_), .B(n253), .C(mem_1__32_), .D(n252), .Z(n254) );
  ND2 U285 ( .A(n255), .B(n254), .Z(rd_data[32]) );
  EO U286 ( .A(wr_ptr[0]), .B(wr_en), .Z(n617) );
  EO U287 ( .A(N45), .B(rd_en), .Z(n421) );
  AO7 U288 ( .A(rd_en), .B(n196), .C(n256), .Z(n420) );
  AO7 U289 ( .A(rd_en), .B(n3), .C(n257), .Z(n419) );
  AO7 U290 ( .A(rd_en), .B(n612), .C(n257), .Z(n418) );
  AO7 U291 ( .A(n615), .B(n256), .C(n258), .Z(n417) );
  MUX21L U292 ( .A(grey_rd_ptr_dly[0]), .B(n259), .S(rd_en), .Z(n258) );
  NR2 U293 ( .A(n260), .B(N45), .Z(n259) );
  AO7 U294 ( .A(rd_en), .B(n611), .C(n261), .Z(n416) );
  IV U295 ( .A(n262), .Z(n261) );
  AO4 U296 ( .A(n263), .B(n256), .C(n257), .D(n260), .Z(n262) );
  ND2 U297 ( .A(rd_en), .B(n263), .Z(n257) );
  ND2 U298 ( .A(rd_en), .B(n260), .Z(n256) );
  EO U299 ( .A(n196), .B(n615), .Z(n260) );
  EN U300 ( .A(n3), .B(n264), .Z(n263) );
  NR2 U301 ( .A(n196), .B(n615), .Z(n264) );
  AO7 U302 ( .A(wr_en), .B(n1), .C(n265), .Z(n415) );
  MUX21L U303 ( .A(n610), .B(n266), .S(n267), .Z(n414) );
  MUX21L U304 ( .A(n609), .B(n268), .S(n267), .Z(n413) );
  MUX21L U305 ( .A(n608), .B(n269), .S(n267), .Z(n412) );
  MUX21L U306 ( .A(n607), .B(n270), .S(n267), .Z(n411) );
  MUX21L U307 ( .A(n606), .B(n271), .S(n267), .Z(n410) );
  MUX21L U308 ( .A(n605), .B(n272), .S(n267), .Z(n409) );
  MUX21L U309 ( .A(n604), .B(n273), .S(n267), .Z(n408) );
  MUX21L U310 ( .A(n603), .B(n274), .S(n267), .Z(n407) );
  MUX21L U311 ( .A(n602), .B(n275), .S(n267), .Z(n406) );
  MUX21L U312 ( .A(n601), .B(n276), .S(n267), .Z(n405) );
  MUX21L U313 ( .A(n600), .B(n277), .S(n267), .Z(n404) );
  MUX21L U314 ( .A(n599), .B(n422), .S(n267), .Z(n403) );
  MUX21L U315 ( .A(n598), .B(n423), .S(n267), .Z(n402) );
  MUX21L U316 ( .A(n597), .B(n424), .S(n267), .Z(n401) );
  MUX21L U317 ( .A(n596), .B(n425), .S(n267), .Z(n400) );
  MUX21L U318 ( .A(n595), .B(n426), .S(n267), .Z(n399) );
  MUX21L U319 ( .A(n594), .B(n427), .S(n267), .Z(n398) );
  MUX21L U320 ( .A(n593), .B(n428), .S(n267), .Z(n397) );
  MUX21L U321 ( .A(n592), .B(n429), .S(n267), .Z(n396) );
  MUX21L U322 ( .A(n591), .B(n430), .S(n267), .Z(n395) );
  MUX21L U323 ( .A(n590), .B(n431), .S(n267), .Z(n394) );
  MUX21L U324 ( .A(n589), .B(n432), .S(n267), .Z(n393) );
  MUX21L U325 ( .A(n588), .B(n433), .S(n267), .Z(n392) );
  MUX21L U326 ( .A(n587), .B(n434), .S(n267), .Z(n391) );
  MUX21L U327 ( .A(n586), .B(n435), .S(n267), .Z(n390) );
  MUX21L U328 ( .A(n585), .B(n436), .S(n267), .Z(n389) );
  MUX21L U329 ( .A(n584), .B(n437), .S(n267), .Z(n388) );
  MUX21L U330 ( .A(n583), .B(n438), .S(n267), .Z(n387) );
  MUX21L U331 ( .A(n582), .B(n439), .S(n267), .Z(n386) );
  MUX21L U332 ( .A(n581), .B(n440), .S(n267), .Z(n385) );
  MUX21L U333 ( .A(n580), .B(n441), .S(n267), .Z(n384) );
  MUX21L U334 ( .A(n579), .B(n442), .S(n267), .Z(n383) );
  MUX21L U335 ( .A(n578), .B(n443), .S(n267), .Z(n382) );
  NR3 U336 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .C(n444), .Z(n267) );
  MUX21L U337 ( .A(n577), .B(n266), .S(n445), .Z(n381) );
  MUX21L U338 ( .A(n576), .B(n268), .S(n445), .Z(n380) );
  MUX21L U339 ( .A(n575), .B(n269), .S(n445), .Z(n379) );
  MUX21L U340 ( .A(n574), .B(n270), .S(n445), .Z(n378) );
  MUX21L U341 ( .A(n573), .B(n271), .S(n445), .Z(n377) );
  MUX21L U342 ( .A(n572), .B(n272), .S(n445), .Z(n376) );
  MUX21L U343 ( .A(n571), .B(n273), .S(n445), .Z(n375) );
  MUX21L U344 ( .A(n570), .B(n274), .S(n445), .Z(n374) );
  MUX21L U345 ( .A(n569), .B(n275), .S(n445), .Z(n373) );
  MUX21L U346 ( .A(n568), .B(n276), .S(n445), .Z(n372) );
  MUX21L U347 ( .A(n567), .B(n277), .S(n445), .Z(n371) );
  MUX21L U348 ( .A(n566), .B(n422), .S(n445), .Z(n370) );
  MUX21L U349 ( .A(n565), .B(n423), .S(n445), .Z(n369) );
  MUX21L U350 ( .A(n564), .B(n424), .S(n445), .Z(n368) );
  MUX21L U351 ( .A(n563), .B(n425), .S(n445), .Z(n367) );
  MUX21L U352 ( .A(n562), .B(n426), .S(n445), .Z(n366) );
  MUX21L U353 ( .A(n561), .B(n427), .S(n445), .Z(n365) );
  MUX21L U354 ( .A(n560), .B(n428), .S(n445), .Z(n364) );
  MUX21L U355 ( .A(n559), .B(n429), .S(n445), .Z(n363) );
  MUX21L U356 ( .A(n558), .B(n430), .S(n445), .Z(n362) );
  MUX21L U357 ( .A(n557), .B(n431), .S(n445), .Z(n361) );
  MUX21L U358 ( .A(n556), .B(n432), .S(n445), .Z(n360) );
  MUX21L U359 ( .A(n555), .B(n433), .S(n445), .Z(n359) );
  MUX21L U360 ( .A(n554), .B(n434), .S(n445), .Z(n358) );
  MUX21L U361 ( .A(n553), .B(n435), .S(n445), .Z(n357) );
  MUX21L U362 ( .A(n552), .B(n436), .S(n445), .Z(n356) );
  MUX21L U363 ( .A(n551), .B(n437), .S(n445), .Z(n355) );
  MUX21L U364 ( .A(n550), .B(n438), .S(n445), .Z(n354) );
  MUX21L U365 ( .A(n549), .B(n439), .S(n445), .Z(n353) );
  MUX21L U366 ( .A(n548), .B(n440), .S(n445), .Z(n352) );
  MUX21L U367 ( .A(n547), .B(n441), .S(n445), .Z(n351) );
  MUX21L U368 ( .A(n546), .B(n442), .S(n445), .Z(n350) );
  MUX21L U369 ( .A(n545), .B(n443), .S(n445), .Z(n349) );
  NR3 U370 ( .A(n4), .B(wr_ptr[1]), .C(n444), .Z(n445) );
  MUX21L U371 ( .A(n544), .B(n266), .S(n446), .Z(n348) );
  MUX21L U372 ( .A(n543), .B(n268), .S(n446), .Z(n347) );
  MUX21L U373 ( .A(n542), .B(n269), .S(n446), .Z(n346) );
  MUX21L U374 ( .A(n541), .B(n270), .S(n446), .Z(n345) );
  MUX21L U375 ( .A(n540), .B(n271), .S(n446), .Z(n344) );
  MUX21L U376 ( .A(n539), .B(n272), .S(n446), .Z(n343) );
  MUX21L U377 ( .A(n538), .B(n273), .S(n446), .Z(n342) );
  MUX21L U378 ( .A(n537), .B(n274), .S(n446), .Z(n341) );
  MUX21L U379 ( .A(n536), .B(n275), .S(n446), .Z(n340) );
  MUX21L U380 ( .A(n535), .B(n276), .S(n446), .Z(n339) );
  MUX21L U381 ( .A(n534), .B(n277), .S(n446), .Z(n338) );
  MUX21L U382 ( .A(n533), .B(n422), .S(n446), .Z(n337) );
  MUX21L U383 ( .A(n532), .B(n423), .S(n446), .Z(n336) );
  MUX21L U384 ( .A(n531), .B(n424), .S(n446), .Z(n335) );
  MUX21L U385 ( .A(n530), .B(n425), .S(n446), .Z(n334) );
  MUX21L U386 ( .A(n529), .B(n426), .S(n446), .Z(n333) );
  MUX21L U387 ( .A(n528), .B(n427), .S(n446), .Z(n332) );
  MUX21L U388 ( .A(n527), .B(n428), .S(n446), .Z(n331) );
  MUX21L U389 ( .A(n526), .B(n429), .S(n446), .Z(n330) );
  MUX21L U390 ( .A(n525), .B(n430), .S(n446), .Z(n329) );
  MUX21L U391 ( .A(n524), .B(n431), .S(n446), .Z(n328) );
  MUX21L U392 ( .A(n523), .B(n432), .S(n446), .Z(n327) );
  MUX21L U393 ( .A(n522), .B(n433), .S(n446), .Z(n326) );
  MUX21L U394 ( .A(n521), .B(n434), .S(n446), .Z(n325) );
  MUX21L U395 ( .A(n520), .B(n435), .S(n446), .Z(n324) );
  MUX21L U396 ( .A(n519), .B(n436), .S(n446), .Z(n323) );
  MUX21L U397 ( .A(n518), .B(n437), .S(n446), .Z(n322) );
  MUX21L U398 ( .A(n517), .B(n438), .S(n446), .Z(n321) );
  MUX21L U399 ( .A(n516), .B(n439), .S(n446), .Z(n320) );
  MUX21L U400 ( .A(n515), .B(n440), .S(n446), .Z(n319) );
  MUX21L U401 ( .A(n514), .B(n441), .S(n446), .Z(n318) );
  MUX21L U402 ( .A(n513), .B(n442), .S(n446), .Z(n317) );
  MUX21L U403 ( .A(n512), .B(n443), .S(n446), .Z(n316) );
  NR3 U404 ( .A(n444), .B(wr_ptr[0]), .C(n1), .Z(n446) );
  MUX21L U405 ( .A(n511), .B(n266), .S(n447), .Z(n315) );
  IV U406 ( .A(wr_data[0]), .Z(n266) );
  MUX21L U407 ( .A(n510), .B(n268), .S(n447), .Z(n314) );
  IV U408 ( .A(wr_data[32]), .Z(n268) );
  MUX21L U409 ( .A(n509), .B(n269), .S(n447), .Z(n313) );
  IV U410 ( .A(wr_data[31]), .Z(n269) );
  MUX21L U411 ( .A(n508), .B(n270), .S(n447), .Z(n312) );
  IV U412 ( .A(wr_data[30]), .Z(n270) );
  MUX21L U413 ( .A(n507), .B(n271), .S(n447), .Z(n311) );
  IV U414 ( .A(wr_data[29]), .Z(n271) );
  MUX21L U415 ( .A(n506), .B(n272), .S(n447), .Z(n310) );
  IV U416 ( .A(wr_data[28]), .Z(n272) );
  MUX21L U417 ( .A(n505), .B(n273), .S(n447), .Z(n309) );
  IV U418 ( .A(wr_data[27]), .Z(n273) );
  MUX21L U419 ( .A(n504), .B(n274), .S(n447), .Z(n308) );
  IV U420 ( .A(wr_data[26]), .Z(n274) );
  MUX21L U421 ( .A(n503), .B(n275), .S(n447), .Z(n307) );
  IV U422 ( .A(wr_data[25]), .Z(n275) );
  MUX21L U423 ( .A(n502), .B(n276), .S(n447), .Z(n306) );
  IV U424 ( .A(wr_data[24]), .Z(n276) );
  MUX21L U425 ( .A(n501), .B(n277), .S(n447), .Z(n305) );
  IV U426 ( .A(wr_data[23]), .Z(n277) );
  MUX21L U427 ( .A(n500), .B(n422), .S(n447), .Z(n304) );
  IV U428 ( .A(wr_data[22]), .Z(n422) );
  MUX21L U429 ( .A(n499), .B(n423), .S(n447), .Z(n303) );
  IV U430 ( .A(wr_data[21]), .Z(n423) );
  MUX21L U431 ( .A(n498), .B(n424), .S(n447), .Z(n302) );
  IV U432 ( .A(wr_data[20]), .Z(n424) );
  MUX21L U433 ( .A(n497), .B(n425), .S(n447), .Z(n301) );
  IV U434 ( .A(wr_data[19]), .Z(n425) );
  MUX21L U435 ( .A(n496), .B(n426), .S(n447), .Z(n300) );
  IV U436 ( .A(wr_data[18]), .Z(n426) );
  MUX21L U437 ( .A(n495), .B(n427), .S(n447), .Z(n299) );
  IV U438 ( .A(wr_data[17]), .Z(n427) );
  MUX21L U439 ( .A(n494), .B(n428), .S(n447), .Z(n298) );
  IV U440 ( .A(wr_data[16]), .Z(n428) );
  MUX21L U441 ( .A(n493), .B(n429), .S(n447), .Z(n297) );
  IV U442 ( .A(wr_data[15]), .Z(n429) );
  MUX21L U443 ( .A(n492), .B(n430), .S(n447), .Z(n296) );
  IV U444 ( .A(wr_data[14]), .Z(n430) );
  MUX21L U445 ( .A(n491), .B(n431), .S(n447), .Z(n295) );
  IV U446 ( .A(wr_data[13]), .Z(n431) );
  MUX21L U447 ( .A(n490), .B(n432), .S(n447), .Z(n294) );
  IV U448 ( .A(wr_data[12]), .Z(n432) );
  MUX21L U449 ( .A(n489), .B(n433), .S(n447), .Z(n293) );
  IV U450 ( .A(wr_data[11]), .Z(n433) );
  MUX21L U451 ( .A(n488), .B(n434), .S(n447), .Z(n292) );
  IV U452 ( .A(wr_data[10]), .Z(n434) );
  MUX21L U453 ( .A(n487), .B(n435), .S(n447), .Z(n291) );
  IV U454 ( .A(wr_data[9]), .Z(n435) );
  MUX21L U455 ( .A(n486), .B(n436), .S(n447), .Z(n290) );
  IV U456 ( .A(wr_data[8]), .Z(n436) );
  MUX21L U457 ( .A(n485), .B(n437), .S(n447), .Z(n289) );
  IV U458 ( .A(wr_data[7]), .Z(n437) );
  MUX21L U459 ( .A(n484), .B(n438), .S(n447), .Z(n288) );
  IV U460 ( .A(wr_data[6]), .Z(n438) );
  MUX21L U461 ( .A(n483), .B(n439), .S(n447), .Z(n287) );
  IV U462 ( .A(wr_data[5]), .Z(n439) );
  MUX21L U463 ( .A(n482), .B(n440), .S(n447), .Z(n286) );
  IV U464 ( .A(wr_data[4]), .Z(n440) );
  MUX21L U465 ( .A(n481), .B(n441), .S(n447), .Z(n285) );
  IV U466 ( .A(wr_data[3]), .Z(n441) );
  MUX21L U467 ( .A(n480), .B(n442), .S(n447), .Z(n284) );
  IV U468 ( .A(wr_data[2]), .Z(n442) );
  MUX21L U469 ( .A(n479), .B(n443), .S(n447), .Z(n283) );
  NR2 U470 ( .A(n448), .B(n444), .Z(n447) );
  IV U471 ( .A(wr_data[1]), .Z(n443) );
  AO7 U472 ( .A(wr_en), .B(n2), .C(n449), .Z(n282) );
  AO7 U473 ( .A(wr_en), .B(n478), .C(n449), .Z(n281) );
  AO7 U474 ( .A(n4), .B(n265), .C(n450), .Z(n280) );
  MUX21L U475 ( .A(grey_wr_ptr[0]), .B(n451), .S(wr_en), .Z(n450) );
  NR2 U476 ( .A(wr_ptr[0]), .B(n452), .Z(n451) );
  AO7 U477 ( .A(test_so5), .B(n265), .C(n453), .Z(n279) );
  EO1 U478 ( .A(grey_wr_ptr[1]), .B(n444), .C(n449), .D(n452), .Z(n453) );
  ND2 U479 ( .A(wr_en), .B(n454), .Z(n449) );
  EN U480 ( .A(test_so5), .B(n448), .Z(n454) );
  ND2 U481 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .Z(n448) );
  ND2 U482 ( .A(wr_en), .B(n452), .Z(n265) );
  EN U483 ( .A(n1), .B(wr_ptr[0]), .Z(n452) );
  AO4 U484 ( .A(n455), .B(n444), .C(n477), .D(n456), .Z(n278) );
  IV U485 ( .A(wr_en), .Z(n444) );
  AN2 U486 ( .A(n457), .B(n477), .Z(n455) );
  AN3 U487 ( .A(n458), .B(n459), .C(n460), .Z(empty) );
  IV U488 ( .A(n461), .Z(n460) );
  IV U489 ( .A(n457), .Z(afull) );
  AO3 U490 ( .A(n462), .B(n463), .C(n464), .D(n456), .Z(n457) );
  EO U491 ( .A(n465), .B(n466), .Z(n456) );
  EN U492 ( .A(sync_rd_ptr_1[2]), .B(n2), .Z(n466) );
  AO5 U493 ( .A(n463), .B(n467), .C(n1), .Z(n465) );
  EO U494 ( .A(sync_rd_ptr_1[2]), .B(sync_rd_ptr_1[1]), .Z(n467) );
  EO U495 ( .A(n468), .B(n469), .Z(n464) );
  EO U496 ( .A(wr_ptr[1]), .B(n463), .Z(n469) );
  NR2 U497 ( .A(wr_ptr[0]), .B(n470), .Z(n463) );
  AN2 U498 ( .A(wr_ptr[0]), .B(n470), .Z(n462) );
  EN U499 ( .A(n468), .B(sync_rd_ptr_1[0]), .Z(n470) );
  EN U500 ( .A(n614), .B(sync_rd_ptr_1[2]), .Z(n468) );
  AN3 U501 ( .A(n459), .B(n461), .C(n458), .Z(aempty) );
  EO U502 ( .A(n471), .B(n472), .Z(n458) );
  NR2 U503 ( .A(n196), .B(n473), .Z(n472) );
  EO U504 ( .A(n3), .B(test_so1), .Z(n471) );
  AO7 U505 ( .A(n474), .B(N45), .C(n473), .Z(n461) );
  EN U506 ( .A(n475), .B(n476), .Z(n459) );
  EO U507 ( .A(n473), .B(n196), .Z(n475) );
  ND2 U508 ( .A(n474), .B(N45), .Z(n473) );
  EN U509 ( .A(n476), .B(sync_wr_ptr_1_0_), .Z(n474) );
  EN U510 ( .A(n616), .B(test_so1), .Z(n476) );
endmodule
