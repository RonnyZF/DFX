module async_fifo_36_8_0_1_test_1 ( wr_clk, wr_reset_n, wr_en, wr_data, full, 
        afull, rd_clk, rd_reset_n, rd_en, empty, aempty, rd_data, test_si8, 
        test_si7, test_si6, test_si5, test_si4, test_si3, test_si2, test_si1, 
        test_so8, test_so7, test_so6, test_so5, test_so4, test_so3, test_so2, 
        test_so1, test_se );
  input [35:0] wr_data;
  output [35:0] rd_data;
  input wr_clk, wr_reset_n, wr_en, rd_clk, rd_reset_n, rd_en, test_si8,
         test_si7, test_si6, test_si5, test_si4, test_si3, test_si2, test_si1,
         test_se;
  output full, afull, empty, aempty, test_so8, test_so7, test_so6, test_so5,
         test_so4, test_so3, test_so2, test_so1;
  wire   N69, N70, N71, wr_ptr_2_, wr_ptr_1_, mem_7__35_, mem_7__34_,
         mem_7__33_, mem_7__32_, mem_7__31_, mem_7__30_, mem_7__29_,
         mem_7__28_, mem_7__27_, mem_7__26_, mem_7__25_, mem_7__24_,
         mem_7__23_, mem_7__22_, mem_7__21_, mem_7__20_, mem_7__19_,
         mem_7__18_, mem_7__17_, mem_7__16_, mem_7__15_, mem_7__14_,
         mem_7__13_, mem_7__12_, mem_7__11_, mem_7__10_, mem_7__9_, mem_7__8_,
         mem_7__7_, mem_7__6_, mem_7__5_, mem_7__4_, mem_7__3_, mem_7__2_,
         mem_7__1_, mem_6__35_, mem_6__34_, mem_6__33_, mem_6__32_, mem_6__31_,
         mem_6__30_, mem_6__29_, mem_6__28_, mem_6__27_, mem_6__26_,
         mem_6__25_, mem_6__24_, mem_6__23_, mem_6__22_, mem_6__21_,
         mem_6__20_, mem_6__19_, mem_6__18_, mem_6__17_, mem_6__16_,
         mem_6__15_, mem_6__14_, mem_6__13_, mem_6__12_, mem_6__11_,
         mem_6__10_, mem_6__9_, mem_6__8_, mem_6__7_, mem_6__6_, mem_6__5_,
         mem_6__4_, mem_6__3_, mem_6__2_, mem_6__1_, mem_6__0_, mem_5__35_,
         mem_5__34_, mem_5__33_, mem_5__32_, mem_5__31_, mem_5__30_,
         mem_5__29_, mem_5__28_, mem_5__27_, mem_5__26_, mem_5__24_,
         mem_5__23_, mem_5__22_, mem_5__21_, mem_5__20_, mem_5__19_,
         mem_5__18_, mem_5__17_, mem_5__16_, mem_5__15_, mem_5__14_,
         mem_5__13_, mem_5__12_, mem_5__11_, mem_5__10_, mem_5__9_, mem_5__8_,
         mem_5__7_, mem_5__6_, mem_5__5_, mem_5__4_, mem_5__3_, mem_5__2_,
         mem_5__1_, mem_5__0_, mem_4__35_, mem_4__34_, mem_4__33_, mem_4__32_,
         mem_4__31_, mem_4__30_, mem_4__29_, mem_4__28_, mem_4__27_,
         mem_4__26_, mem_4__25_, mem_4__24_, mem_4__23_, mem_4__22_,
         mem_4__21_, mem_4__20_, mem_4__19_, mem_4__18_, mem_4__17_,
         mem_4__16_, mem_4__15_, mem_4__13_, mem_4__12_, mem_4__11_,
         mem_4__10_, mem_4__9_, mem_4__8_, mem_4__7_, mem_4__6_, mem_4__5_,
         mem_4__4_, mem_4__3_, mem_4__2_, mem_4__1_, mem_4__0_, mem_3__35_,
         mem_3__34_, mem_3__33_, mem_3__32_, mem_3__31_, mem_3__30_,
         mem_3__29_, mem_3__28_, mem_3__27_, mem_3__26_, mem_3__25_,
         mem_3__24_, mem_3__23_, mem_3__22_, mem_3__21_, mem_3__20_,
         mem_3__19_, mem_3__18_, mem_3__17_, mem_3__16_, mem_3__15_,
         mem_3__14_, mem_3__13_, mem_3__12_, mem_3__11_, mem_3__10_, mem_3__9_,
         mem_3__8_, mem_3__7_, mem_3__6_, mem_3__5_, mem_3__4_, mem_3__2_,
         mem_3__1_, mem_3__0_, mem_2__35_, mem_2__34_, mem_2__33_, mem_2__32_,
         mem_2__31_, mem_2__30_, mem_2__29_, mem_2__28_, mem_2__27_,
         mem_2__26_, mem_2__25_, mem_2__24_, mem_2__23_, mem_2__22_,
         mem_2__21_, mem_2__20_, mem_2__19_, mem_2__18_, mem_2__17_,
         mem_2__16_, mem_2__15_, mem_2__14_, mem_2__13_, mem_2__12_,
         mem_2__11_, mem_2__10_, mem_2__9_, mem_2__8_, mem_2__7_, mem_2__6_,
         mem_2__5_, mem_2__4_, mem_2__3_, mem_2__2_, mem_2__1_, mem_2__0_,
         mem_1__35_, mem_1__34_, mem_1__33_, mem_1__32_, mem_1__31_,
         mem_1__30_, mem_1__29_, mem_1__27_, mem_1__26_, mem_1__25_,
         mem_1__24_, mem_1__23_, mem_1__22_, mem_1__21_, mem_1__20_,
         mem_1__19_, mem_1__18_, mem_1__17_, mem_1__16_, mem_1__15_,
         mem_1__14_, mem_1__13_, mem_1__12_, mem_1__11_, mem_1__10_, mem_1__9_,
         mem_1__8_, mem_1__7_, mem_1__6_, mem_1__5_, mem_1__4_, mem_1__3_,
         mem_1__2_, mem_1__1_, mem_1__0_, mem_0__35_, mem_0__34_, mem_0__33_,
         mem_0__32_, mem_0__31_, mem_0__30_, mem_0__29_, mem_0__28_,
         mem_0__27_, mem_0__26_, mem_0__25_, mem_0__24_, mem_0__23_,
         mem_0__22_, mem_0__21_, mem_0__20_, mem_0__19_, mem_0__18_,
         mem_0__17_, mem_0__15_, mem_0__14_, mem_0__13_, mem_0__12_,
         mem_0__11_, mem_0__10_, mem_0__9_, mem_0__8_, mem_0__7_, mem_0__6_,
         mem_0__5_, mem_0__4_, mem_0__3_, mem_0__2_, mem_0__1_, mem_0__0_,
         rd_ptr_3_1, sync_wr_ptr_1_1_, sync_wr_ptr_1_0_, n360, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n356,
         n357, n358, n359, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1244;
  wire   [3:0] grey_wr_ptr;
  wire   [3:0] grey_rd_ptr_dly;
  wire   [3:0] sync_rd_ptr_1;
  wire   [3:0] sync_rd_ptr_0;
  wire   [3:0] sync_wr_ptr_0;

  FD2S sync_wr_ptr_1_reg_2_ ( .D(sync_wr_ptr_0[2]), .TI(sync_wr_ptr_1_1_), 
        .TE(test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(n1244), .QN(n971) );
  FD1S mem_reg_7__35_ ( .D(n498), .TI(mem_7__34_), .TE(test_se), .CP(n15), .Q(
        mem_7__35_), .QN(n1012) );
  FD1S mem_reg_7__34_ ( .D(n497), .TI(mem_7__33_), .TE(test_se), .CP(n15), .Q(
        mem_7__34_), .QN(n1011) );
  FD1S mem_reg_7__33_ ( .D(n496), .TI(mem_7__32_), .TE(test_se), .CP(n14), .Q(
        mem_7__33_), .QN(n1010) );
  FD1S mem_reg_7__32_ ( .D(n495), .TI(mem_7__31_), .TE(test_se), .CP(n14), .Q(
        mem_7__32_), .QN(n1009) );
  FD1S mem_reg_7__31_ ( .D(n494), .TI(mem_7__30_), .TE(test_se), .CP(n14), .Q(
        mem_7__31_), .QN(n1008) );
  FD1S mem_reg_7__30_ ( .D(n493), .TI(mem_7__29_), .TE(test_se), .CP(n14), .Q(
        mem_7__30_), .QN(n1007) );
  FD1S mem_reg_7__29_ ( .D(n492), .TI(mem_7__28_), .TE(test_se), .CP(n14), .Q(
        mem_7__29_), .QN(n1006) );
  FD1S mem_reg_7__28_ ( .D(n491), .TI(mem_7__27_), .TE(test_se), .CP(n14), .Q(
        mem_7__28_), .QN(n1005) );
  FD1S mem_reg_7__27_ ( .D(n490), .TI(mem_7__26_), .TE(test_se), .CP(n14), .Q(
        mem_7__27_), .QN(n1004) );
  FD1S mem_reg_7__26_ ( .D(n489), .TI(mem_7__25_), .TE(test_se), .CP(n14), .Q(
        mem_7__26_), .QN(n1003) );
  FD1S mem_reg_7__25_ ( .D(n488), .TI(mem_7__24_), .TE(test_se), .CP(n14), .Q(
        mem_7__25_), .QN(n1002) );
  FD1S mem_reg_7__24_ ( .D(n487), .TI(mem_7__23_), .TE(test_se), .CP(n14), .Q(
        mem_7__24_), .QN(n1001) );
  FD1S mem_reg_7__23_ ( .D(n486), .TI(mem_7__22_), .TE(test_se), .CP(n14), .Q(
        mem_7__23_), .QN(n1000) );
  FD1S mem_reg_7__22_ ( .D(n485), .TI(mem_7__21_), .TE(test_se), .CP(n14), .Q(
        mem_7__22_), .QN(n999) );
  FD1S mem_reg_7__21_ ( .D(n484), .TI(mem_7__20_), .TE(test_se), .CP(n13), .Q(
        mem_7__21_), .QN(n998) );
  FD1S mem_reg_7__20_ ( .D(n483), .TI(mem_7__19_), .TE(test_se), .CP(n13), .Q(
        mem_7__20_), .QN(n997) );
  FD1S mem_reg_7__19_ ( .D(n482), .TI(mem_7__18_), .TE(test_se), .CP(n13), .Q(
        mem_7__19_), .QN(n996) );
  FD1S mem_reg_7__18_ ( .D(n481), .TI(mem_7__17_), .TE(test_se), .CP(n13), .Q(
        mem_7__18_), .QN(n995) );
  FD1S mem_reg_7__17_ ( .D(n480), .TI(mem_7__16_), .TE(test_se), .CP(n13), .Q(
        mem_7__17_), .QN(n994) );
  FD1S mem_reg_7__16_ ( .D(n479), .TI(mem_7__15_), .TE(test_se), .CP(n13), .Q(
        mem_7__16_), .QN(n993) );
  FD1S mem_reg_7__15_ ( .D(n478), .TI(mem_7__14_), .TE(test_se), .CP(n13), .Q(
        mem_7__15_), .QN(n992) );
  FD1S mem_reg_7__14_ ( .D(n477), .TI(mem_7__13_), .TE(test_se), .CP(n13), .Q(
        mem_7__14_), .QN(n991) );
  FD1S mem_reg_7__13_ ( .D(n476), .TI(mem_7__12_), .TE(test_se), .CP(n13), .Q(
        mem_7__13_), .QN(n990) );
  FD1S mem_reg_7__12_ ( .D(n475), .TI(mem_7__11_), .TE(test_se), .CP(n13), .Q(
        mem_7__12_), .QN(n989) );
  FD1S mem_reg_7__11_ ( .D(n474), .TI(mem_7__10_), .TE(test_se), .CP(n13), .Q(
        mem_7__11_), .QN(n988) );
  FD1S mem_reg_7__10_ ( .D(n473), .TI(mem_7__9_), .TE(test_se), .CP(n13), .Q(
        mem_7__10_), .QN(n987) );
  FD1S mem_reg_7__9_ ( .D(n472), .TI(mem_7__8_), .TE(test_se), .CP(n12), .Q(
        mem_7__9_), .QN(n986) );
  FD1S mem_reg_7__8_ ( .D(n471), .TI(mem_7__7_), .TE(test_se), .CP(n12), .Q(
        mem_7__8_), .QN(n985) );
  FD1S mem_reg_7__7_ ( .D(n470), .TI(mem_7__6_), .TE(test_se), .CP(n12), .Q(
        mem_7__7_), .QN(n984) );
  FD1S mem_reg_7__6_ ( .D(n469), .TI(mem_7__5_), .TE(test_se), .CP(n12), .Q(
        mem_7__6_), .QN(n983) );
  FD1S mem_reg_7__5_ ( .D(n468), .TI(mem_7__4_), .TE(test_se), .CP(n12), .Q(
        mem_7__5_), .QN(n982) );
  FD1S mem_reg_7__4_ ( .D(n467), .TI(mem_7__3_), .TE(test_se), .CP(n12), .Q(
        mem_7__4_), .QN(n981) );
  FD1S mem_reg_7__3_ ( .D(n466), .TI(mem_7__2_), .TE(test_se), .CP(n12), .Q(
        mem_7__3_), .QN(n980) );
  FD1S mem_reg_7__2_ ( .D(n465), .TI(mem_7__1_), .TE(test_se), .CP(n12), .Q(
        mem_7__2_), .QN(n979) );
  FD1S mem_reg_7__1_ ( .D(n464), .TI(test_si7), .TE(test_se), .CP(n12), .Q(
        mem_7__1_), .QN(n978) );
  FD1S mem_reg_7__0_ ( .D(n499), .TI(mem_6__35_), .TE(test_se), .CP(n15), .Q(
        test_so6), .QN(n1013) );
  FD1S mem_reg_6__35_ ( .D(n534), .TI(mem_6__34_), .TE(test_se), .CP(n11), .Q(
        mem_6__35_), .QN(n1048) );
  FD1S mem_reg_6__34_ ( .D(n533), .TI(mem_6__33_), .TE(test_se), .CP(n11), .Q(
        mem_6__34_), .QN(n1047) );
  FD1S mem_reg_6__33_ ( .D(n532), .TI(mem_6__32_), .TE(test_se), .CP(n11), .Q(
        mem_6__33_), .QN(n1046) );
  FD1S mem_reg_6__32_ ( .D(n531), .TI(mem_6__31_), .TE(test_se), .CP(n11), .Q(
        mem_6__32_), .QN(n1045) );
  FD1S mem_reg_6__31_ ( .D(n530), .TI(mem_6__30_), .TE(test_se), .CP(n11), .Q(
        mem_6__31_), .QN(n1044) );
  FD1S mem_reg_6__30_ ( .D(n529), .TI(mem_6__29_), .TE(test_se), .CP(n11), .Q(
        mem_6__30_), .QN(n1043) );
  FD1S mem_reg_6__29_ ( .D(n528), .TI(mem_6__28_), .TE(test_se), .CP(n11), .Q(
        mem_6__29_), .QN(n1042) );
  FD1S mem_reg_6__28_ ( .D(n527), .TI(mem_6__27_), .TE(test_se), .CP(n11), .Q(
        mem_6__28_), .QN(n1041) );
  FD1S mem_reg_6__27_ ( .D(n526), .TI(mem_6__26_), .TE(test_se), .CP(n11), .Q(
        mem_6__27_), .QN(n1040) );
  FD1S mem_reg_6__26_ ( .D(n525), .TI(mem_6__25_), .TE(test_se), .CP(n11), .Q(
        mem_6__26_), .QN(n1039) );
  FD1S mem_reg_6__25_ ( .D(n524), .TI(mem_6__24_), .TE(test_se), .CP(n11), .Q(
        mem_6__25_), .QN(n1038) );
  FD1S mem_reg_6__24_ ( .D(n523), .TI(mem_6__23_), .TE(test_se), .CP(n11), .Q(
        mem_6__24_), .QN(n1037) );
  FD1S mem_reg_6__23_ ( .D(n522), .TI(mem_6__22_), .TE(test_se), .CP(n10), .Q(
        mem_6__23_), .QN(n1036) );
  FD1S mem_reg_6__22_ ( .D(n521), .TI(mem_6__21_), .TE(test_se), .CP(n10), .Q(
        mem_6__22_), .QN(n1035) );
  FD1S mem_reg_6__21_ ( .D(n520), .TI(mem_6__20_), .TE(test_se), .CP(n10), .Q(
        mem_6__21_), .QN(n1034) );
  FD1S mem_reg_6__20_ ( .D(n519), .TI(mem_6__19_), .TE(test_se), .CP(n10), .Q(
        mem_6__20_), .QN(n1033) );
  FD1S mem_reg_6__19_ ( .D(n518), .TI(mem_6__18_), .TE(test_se), .CP(n10), .Q(
        mem_6__19_), .QN(n1032) );
  FD1S mem_reg_6__18_ ( .D(n517), .TI(mem_6__17_), .TE(test_se), .CP(n10), .Q(
        mem_6__18_), .QN(n1031) );
  FD1S mem_reg_6__17_ ( .D(n516), .TI(mem_6__16_), .TE(test_se), .CP(n10), .Q(
        mem_6__17_), .QN(n1030) );
  FD1S mem_reg_6__16_ ( .D(n515), .TI(mem_6__15_), .TE(test_se), .CP(n10), .Q(
        mem_6__16_), .QN(n1029) );
  FD1S mem_reg_6__15_ ( .D(n514), .TI(mem_6__14_), .TE(test_se), .CP(n10), .Q(
        mem_6__15_), .QN(n1028) );
  FD1S mem_reg_6__14_ ( .D(n513), .TI(mem_6__13_), .TE(test_se), .CP(n10), .Q(
        mem_6__14_), .QN(n1027) );
  FD1S mem_reg_6__13_ ( .D(n512), .TI(mem_6__12_), .TE(test_se), .CP(n10), .Q(
        mem_6__13_), .QN(n1026) );
  FD1S mem_reg_6__12_ ( .D(n511), .TI(mem_6__11_), .TE(test_se), .CP(n10), .Q(
        mem_6__12_), .QN(n1025) );
  FD1S mem_reg_6__11_ ( .D(n510), .TI(mem_6__10_), .TE(test_se), .CP(n9), .Q(
        mem_6__11_), .QN(n1024) );
  FD1S mem_reg_6__10_ ( .D(n509), .TI(mem_6__9_), .TE(test_se), .CP(n9), .Q(
        mem_6__10_), .QN(n1023) );
  FD1S mem_reg_6__9_ ( .D(n508), .TI(mem_6__8_), .TE(test_se), .CP(n9), .Q(
        mem_6__9_), .QN(n1022) );
  FD1S mem_reg_6__8_ ( .D(n507), .TI(mem_6__7_), .TE(test_se), .CP(n9), .Q(
        mem_6__8_), .QN(n1021) );
  FD1S mem_reg_6__7_ ( .D(n506), .TI(mem_6__6_), .TE(test_se), .CP(n9), .Q(
        mem_6__7_), .QN(n1020) );
  FD1S mem_reg_6__6_ ( .D(n505), .TI(mem_6__5_), .TE(test_se), .CP(n9), .Q(
        mem_6__6_), .QN(n1019) );
  FD1S mem_reg_6__5_ ( .D(n504), .TI(mem_6__4_), .TE(test_se), .CP(n9), .Q(
        mem_6__5_), .QN(n1018) );
  FD1S mem_reg_6__4_ ( .D(n503), .TI(mem_6__3_), .TE(test_se), .CP(n9), .Q(
        mem_6__4_), .QN(n1017) );
  FD1S mem_reg_6__3_ ( .D(n502), .TI(mem_6__2_), .TE(test_se), .CP(n9), .Q(
        mem_6__3_), .QN(n1016) );
  FD1S mem_reg_6__2_ ( .D(n501), .TI(mem_6__1_), .TE(test_se), .CP(n9), .Q(
        mem_6__2_), .QN(n1015) );
  FD1S mem_reg_6__1_ ( .D(n500), .TI(mem_6__0_), .TE(test_se), .CP(n9), .Q(
        mem_6__1_), .QN(n1014) );
  FD1S mem_reg_6__0_ ( .D(n535), .TI(mem_5__35_), .TE(test_se), .CP(n12), .Q(
        mem_6__0_), .QN(n1049) );
  FD1S mem_reg_5__35_ ( .D(n570), .TI(mem_5__34_), .TE(test_se), .CP(n8), .Q(
        mem_5__35_), .QN(n1084) );
  FD1S mem_reg_5__34_ ( .D(n569), .TI(mem_5__33_), .TE(test_se), .CP(n8), .Q(
        mem_5__34_), .QN(n1083) );
  FD1S mem_reg_5__33_ ( .D(n568), .TI(mem_5__32_), .TE(test_se), .CP(n8), .Q(
        mem_5__33_), .QN(n1082) );
  FD1S mem_reg_5__32_ ( .D(n567), .TI(mem_5__31_), .TE(test_se), .CP(n8), .Q(
        mem_5__32_), .QN(n1081) );
  FD1S mem_reg_5__31_ ( .D(n566), .TI(mem_5__30_), .TE(test_se), .CP(n8), .Q(
        mem_5__31_), .QN(n1080) );
  FD1S mem_reg_5__30_ ( .D(n565), .TI(mem_5__29_), .TE(test_se), .CP(n8), .Q(
        mem_5__30_), .QN(n1079) );
  FD1S mem_reg_5__29_ ( .D(n564), .TI(mem_5__28_), .TE(test_se), .CP(n8), .Q(
        mem_5__29_), .QN(n1078) );
  FD1S mem_reg_5__28_ ( .D(n563), .TI(mem_5__27_), .TE(test_se), .CP(n8), .Q(
        mem_5__28_), .QN(n1077) );
  FD1S mem_reg_5__27_ ( .D(n562), .TI(mem_5__26_), .TE(test_se), .CP(n8), .Q(
        mem_5__27_), .QN(n1076) );
  FD1S mem_reg_5__26_ ( .D(n561), .TI(test_si6), .TE(test_se), .CP(n8), .Q(
        mem_5__26_), .QN(n1075) );
  FD1S mem_reg_5__25_ ( .D(n560), .TI(mem_5__24_), .TE(test_se), .CP(n8), .Q(
        test_so5), .QN(n1074) );
  FD1S mem_reg_5__24_ ( .D(n559), .TI(mem_5__23_), .TE(test_se), .CP(n8), .Q(
        mem_5__24_), .QN(n1073) );
  FD1S mem_reg_5__23_ ( .D(n558), .TI(mem_5__22_), .TE(test_se), .CP(n7), .Q(
        mem_5__23_), .QN(n1072) );
  FD1S mem_reg_5__22_ ( .D(n557), .TI(mem_5__21_), .TE(test_se), .CP(n7), .Q(
        mem_5__22_), .QN(n1071) );
  FD1S mem_reg_5__21_ ( .D(n556), .TI(mem_5__20_), .TE(test_se), .CP(n7), .Q(
        mem_5__21_), .QN(n1070) );
  FD1S mem_reg_5__20_ ( .D(n555), .TI(mem_5__19_), .TE(test_se), .CP(n7), .Q(
        mem_5__20_), .QN(n1069) );
  FD1S mem_reg_5__19_ ( .D(n554), .TI(mem_5__18_), .TE(test_se), .CP(n7), .Q(
        mem_5__19_), .QN(n1068) );
  FD1S mem_reg_5__18_ ( .D(n553), .TI(mem_5__17_), .TE(test_se), .CP(n7), .Q(
        mem_5__18_), .QN(n1067) );
  FD1S mem_reg_5__17_ ( .D(n552), .TI(mem_5__16_), .TE(test_se), .CP(n7), .Q(
        mem_5__17_), .QN(n1066) );
  FD1S mem_reg_5__16_ ( .D(n551), .TI(mem_5__15_), .TE(test_se), .CP(n7), .Q(
        mem_5__16_), .QN(n1065) );
  FD1S mem_reg_5__15_ ( .D(n550), .TI(mem_5__14_), .TE(test_se), .CP(n7), .Q(
        mem_5__15_), .QN(n1064) );
  FD1S mem_reg_5__14_ ( .D(n549), .TI(mem_5__13_), .TE(test_se), .CP(n7), .Q(
        mem_5__14_), .QN(n1063) );
  FD1S mem_reg_5__13_ ( .D(n548), .TI(mem_5__12_), .TE(test_se), .CP(n7), .Q(
        mem_5__13_), .QN(n1062) );
  FD1S mem_reg_5__12_ ( .D(n547), .TI(mem_5__11_), .TE(test_se), .CP(n7), .Q(
        mem_5__12_), .QN(n1061) );
  FD1S mem_reg_5__11_ ( .D(n546), .TI(mem_5__10_), .TE(test_se), .CP(n6), .Q(
        mem_5__11_), .QN(n1060) );
  FD1S mem_reg_5__10_ ( .D(n545), .TI(mem_5__9_), .TE(test_se), .CP(n6), .Q(
        mem_5__10_), .QN(n1059) );
  FD1S mem_reg_5__9_ ( .D(n544), .TI(mem_5__8_), .TE(test_se), .CP(n6), .Q(
        mem_5__9_), .QN(n1058) );
  FD1S mem_reg_5__8_ ( .D(n543), .TI(mem_5__7_), .TE(test_se), .CP(n6), .Q(
        mem_5__8_), .QN(n1057) );
  FD1S mem_reg_5__7_ ( .D(n542), .TI(mem_5__6_), .TE(test_se), .CP(n6), .Q(
        mem_5__7_), .QN(n1056) );
  FD1S mem_reg_5__6_ ( .D(n541), .TI(mem_5__5_), .TE(test_se), .CP(n6), .Q(
        mem_5__6_), .QN(n1055) );
  FD1S mem_reg_5__5_ ( .D(n540), .TI(mem_5__4_), .TE(test_se), .CP(n6), .Q(
        mem_5__5_), .QN(n1054) );
  FD1S mem_reg_5__4_ ( .D(n539), .TI(mem_5__3_), .TE(test_se), .CP(n6), .Q(
        mem_5__4_), .QN(n1053) );
  FD1S mem_reg_5__3_ ( .D(n538), .TI(mem_5__2_), .TE(test_se), .CP(n6), .Q(
        mem_5__3_), .QN(n1052) );
  FD1S mem_reg_5__2_ ( .D(n537), .TI(mem_5__1_), .TE(test_se), .CP(n6), .Q(
        mem_5__2_), .QN(n1051) );
  FD1S mem_reg_5__1_ ( .D(n536), .TI(mem_5__0_), .TE(test_se), .CP(n6), .Q(
        mem_5__1_), .QN(n1050) );
  FD1S mem_reg_5__0_ ( .D(n571), .TI(mem_4__35_), .TE(test_se), .CP(n9), .Q(
        mem_5__0_), .QN(n1085) );
  FD1S mem_reg_4__35_ ( .D(n606), .TI(mem_4__34_), .TE(test_se), .CP(n27), .Q(
        mem_4__35_), .QN(n1120) );
  FD1S mem_reg_4__34_ ( .D(n605), .TI(mem_4__33_), .TE(test_se), .CP(n27), .Q(
        mem_4__34_), .QN(n1119) );
  FD1S mem_reg_4__33_ ( .D(n604), .TI(mem_4__32_), .TE(test_se), .CP(n27), .Q(
        mem_4__33_), .QN(n1118) );
  FD1S mem_reg_4__32_ ( .D(n603), .TI(mem_4__31_), .TE(test_se), .CP(n27), .Q(
        mem_4__32_), .QN(n1117) );
  FD1S mem_reg_4__31_ ( .D(n602), .TI(mem_4__30_), .TE(test_se), .CP(n26), .Q(
        mem_4__31_), .QN(n1116) );
  FD1S mem_reg_4__30_ ( .D(n601), .TI(mem_4__29_), .TE(test_se), .CP(n26), .Q(
        mem_4__30_), .QN(n1115) );
  FD1S mem_reg_4__29_ ( .D(n600), .TI(mem_4__28_), .TE(test_se), .CP(n26), .Q(
        mem_4__29_), .QN(n1114) );
  FD1S mem_reg_4__28_ ( .D(n599), .TI(mem_4__27_), .TE(test_se), .CP(n26), .Q(
        mem_4__28_), .QN(n1113) );
  FD1S mem_reg_4__27_ ( .D(n598), .TI(mem_4__26_), .TE(test_se), .CP(n26), .Q(
        mem_4__27_), .QN(n1112) );
  FD1S mem_reg_4__26_ ( .D(n597), .TI(mem_4__25_), .TE(test_se), .CP(n26), .Q(
        mem_4__26_), .QN(n1111) );
  FD1S mem_reg_4__25_ ( .D(n596), .TI(mem_4__24_), .TE(test_se), .CP(n26), .Q(
        mem_4__25_), .QN(n1110) );
  FD1S mem_reg_4__24_ ( .D(n595), .TI(mem_4__23_), .TE(test_se), .CP(n26), .Q(
        mem_4__24_), .QN(n1109) );
  FD1S mem_reg_4__23_ ( .D(n594), .TI(mem_4__22_), .TE(test_se), .CP(n26), .Q(
        mem_4__23_), .QN(n1108) );
  FD1S mem_reg_4__22_ ( .D(n593), .TI(mem_4__21_), .TE(test_se), .CP(n26), .Q(
        mem_4__22_), .QN(n1107) );
  FD1S mem_reg_4__21_ ( .D(n592), .TI(mem_4__20_), .TE(test_se), .CP(n26), .Q(
        mem_4__21_), .QN(n1106) );
  FD1S mem_reg_4__20_ ( .D(n591), .TI(mem_4__19_), .TE(test_se), .CP(n26), .Q(
        mem_4__20_), .QN(n1105) );
  FD1S mem_reg_4__19_ ( .D(n590), .TI(mem_4__18_), .TE(test_se), .CP(n25), .Q(
        mem_4__19_), .QN(n1104) );
  FD1S mem_reg_4__18_ ( .D(n589), .TI(mem_4__17_), .TE(test_se), .CP(n25), .Q(
        mem_4__18_), .QN(n1103) );
  FD1S mem_reg_4__17_ ( .D(n588), .TI(mem_4__16_), .TE(test_se), .CP(n25), .Q(
        mem_4__17_), .QN(n1102) );
  FD1S mem_reg_4__16_ ( .D(n587), .TI(mem_4__15_), .TE(test_se), .CP(n25), .Q(
        mem_4__16_), .QN(n1101) );
  FD1S mem_reg_4__15_ ( .D(n586), .TI(test_si5), .TE(test_se), .CP(n25), .Q(
        mem_4__15_), .QN(n1100) );
  FD1S mem_reg_4__14_ ( .D(n585), .TI(mem_4__13_), .TE(test_se), .CP(n25), .Q(
        test_so4), .QN(n1099) );
  FD1S mem_reg_4__13_ ( .D(n584), .TI(mem_4__12_), .TE(test_se), .CP(n25), .Q(
        mem_4__13_), .QN(n1098) );
  FD1S mem_reg_4__12_ ( .D(n583), .TI(mem_4__11_), .TE(test_se), .CP(n25), .Q(
        mem_4__12_), .QN(n1097) );
  FD1S mem_reg_4__11_ ( .D(n582), .TI(mem_4__10_), .TE(test_se), .CP(n25), .Q(
        mem_4__11_), .QN(n1096) );
  FD1S mem_reg_4__10_ ( .D(n581), .TI(mem_4__9_), .TE(test_se), .CP(n25), .Q(
        mem_4__10_), .QN(n1095) );
  FD1S mem_reg_4__9_ ( .D(n580), .TI(mem_4__8_), .TE(test_se), .CP(n25), .Q(
        mem_4__9_), .QN(n1094) );
  FD1S mem_reg_4__8_ ( .D(n579), .TI(mem_4__7_), .TE(test_se), .CP(n25), .Q(
        mem_4__8_), .QN(n1093) );
  FD1S mem_reg_4__7_ ( .D(n578), .TI(mem_4__6_), .TE(test_se), .CP(n24), .Q(
        mem_4__7_), .QN(n1092) );
  FD1S mem_reg_4__6_ ( .D(n577), .TI(mem_4__5_), .TE(test_se), .CP(n24), .Q(
        mem_4__6_), .QN(n1091) );
  FD1S mem_reg_4__5_ ( .D(n576), .TI(mem_4__4_), .TE(test_se), .CP(n24), .Q(
        mem_4__5_), .QN(n1090) );
  FD1S mem_reg_4__4_ ( .D(n575), .TI(mem_4__3_), .TE(test_se), .CP(n24), .Q(
        mem_4__4_), .QN(n1089) );
  FD1S mem_reg_4__3_ ( .D(n574), .TI(mem_4__2_), .TE(test_se), .CP(n24), .Q(
        mem_4__3_), .QN(n1088) );
  FD1S mem_reg_4__2_ ( .D(n573), .TI(mem_4__1_), .TE(test_se), .CP(n24), .Q(
        mem_4__2_), .QN(n1087) );
  FD1S mem_reg_4__1_ ( .D(n572), .TI(mem_4__0_), .TE(test_se), .CP(n24), .Q(
        mem_4__1_), .QN(n1086) );
  FD1S mem_reg_4__0_ ( .D(n607), .TI(mem_3__35_), .TE(test_se), .CP(n27), .Q(
        mem_4__0_), .QN(n1121) );
  FD1S mem_reg_3__35_ ( .D(n642), .TI(mem_3__34_), .TE(test_se), .CP(n24), .Q(
        mem_3__35_), .QN(n1156) );
  FD1S mem_reg_3__34_ ( .D(n641), .TI(mem_3__33_), .TE(test_se), .CP(n24), .Q(
        mem_3__34_), .QN(n1155) );
  FD1S mem_reg_3__33_ ( .D(n640), .TI(mem_3__32_), .TE(test_se), .CP(n24), .Q(
        mem_3__33_), .QN(n1154) );
  FD1S mem_reg_3__32_ ( .D(n639), .TI(mem_3__31_), .TE(test_se), .CP(n24), .Q(
        mem_3__32_), .QN(n1153) );
  FD1S mem_reg_3__31_ ( .D(n638), .TI(mem_3__30_), .TE(test_se), .CP(n23), .Q(
        mem_3__31_), .QN(n1152) );
  FD1S mem_reg_3__30_ ( .D(n637), .TI(mem_3__29_), .TE(test_se), .CP(n23), .Q(
        mem_3__30_), .QN(n1151) );
  FD1S mem_reg_3__29_ ( .D(n636), .TI(mem_3__28_), .TE(test_se), .CP(n23), .Q(
        mem_3__29_), .QN(n1150) );
  FD1S mem_reg_3__28_ ( .D(n635), .TI(mem_3__27_), .TE(test_se), .CP(n23), .Q(
        mem_3__28_), .QN(n1149) );
  FD1S mem_reg_3__27_ ( .D(n634), .TI(mem_3__26_), .TE(test_se), .CP(n23), .Q(
        mem_3__27_), .QN(n1148) );
  FD1S mem_reg_3__26_ ( .D(n633), .TI(mem_3__25_), .TE(test_se), .CP(n23), .Q(
        mem_3__26_), .QN(n1147) );
  FD1S mem_reg_3__25_ ( .D(n632), .TI(mem_3__24_), .TE(test_se), .CP(n23), .Q(
        mem_3__25_), .QN(n1146) );
  FD1S mem_reg_3__24_ ( .D(n631), .TI(mem_3__23_), .TE(test_se), .CP(n23), .Q(
        mem_3__24_), .QN(n1145) );
  FD1S mem_reg_3__23_ ( .D(n630), .TI(mem_3__22_), .TE(test_se), .CP(n23), .Q(
        mem_3__23_), .QN(n1144) );
  FD1S mem_reg_3__22_ ( .D(n629), .TI(mem_3__21_), .TE(test_se), .CP(n23), .Q(
        mem_3__22_), .QN(n1143) );
  FD1S mem_reg_3__21_ ( .D(n628), .TI(mem_3__20_), .TE(test_se), .CP(n23), .Q(
        mem_3__21_), .QN(n1142) );
  FD1S mem_reg_3__20_ ( .D(n627), .TI(mem_3__19_), .TE(test_se), .CP(n23), .Q(
        mem_3__20_), .QN(n1141) );
  FD1S mem_reg_3__19_ ( .D(n626), .TI(mem_3__18_), .TE(test_se), .CP(n22), .Q(
        mem_3__19_), .QN(n1140) );
  FD1S mem_reg_3__18_ ( .D(n625), .TI(mem_3__17_), .TE(test_se), .CP(n22), .Q(
        mem_3__18_), .QN(n1139) );
  FD1S mem_reg_3__17_ ( .D(n624), .TI(mem_3__16_), .TE(test_se), .CP(n22), .Q(
        mem_3__17_), .QN(n1138) );
  FD1S mem_reg_3__16_ ( .D(n623), .TI(mem_3__15_), .TE(test_se), .CP(n22), .Q(
        mem_3__16_), .QN(n1137) );
  FD1S mem_reg_3__15_ ( .D(n622), .TI(mem_3__14_), .TE(test_se), .CP(n22), .Q(
        mem_3__15_), .QN(n1136) );
  FD1S mem_reg_3__14_ ( .D(n621), .TI(mem_3__13_), .TE(test_se), .CP(n22), .Q(
        mem_3__14_), .QN(n1135) );
  FD1S mem_reg_3__13_ ( .D(n620), .TI(mem_3__12_), .TE(test_se), .CP(n22), .Q(
        mem_3__13_), .QN(n1134) );
  FD1S mem_reg_3__12_ ( .D(n619), .TI(mem_3__11_), .TE(test_se), .CP(n22), .Q(
        mem_3__12_), .QN(n1133) );
  FD1S mem_reg_3__11_ ( .D(n618), .TI(mem_3__10_), .TE(test_se), .CP(n22), .Q(
        mem_3__11_), .QN(n1132) );
  FD1S mem_reg_3__10_ ( .D(n617), .TI(mem_3__9_), .TE(test_se), .CP(n22), .Q(
        mem_3__10_), .QN(n1131) );
  FD1S mem_reg_3__9_ ( .D(n616), .TI(mem_3__8_), .TE(test_se), .CP(n22), .Q(
        mem_3__9_), .QN(n1130) );
  FD1S mem_reg_3__8_ ( .D(n615), .TI(mem_3__7_), .TE(test_se), .CP(n22), .Q(
        mem_3__8_), .QN(n1129) );
  FD1S mem_reg_3__7_ ( .D(n614), .TI(mem_3__6_), .TE(test_se), .CP(n21), .Q(
        mem_3__7_), .QN(n1128) );
  FD1S mem_reg_3__6_ ( .D(n613), .TI(mem_3__5_), .TE(test_se), .CP(n21), .Q(
        mem_3__6_), .QN(n1127) );
  FD1S mem_reg_3__5_ ( .D(n612), .TI(mem_3__4_), .TE(test_se), .CP(n21), .Q(
        mem_3__5_), .QN(n1126) );
  FD1S mem_reg_3__4_ ( .D(n611), .TI(test_si4), .TE(test_se), .CP(n21), .Q(
        mem_3__4_), .QN(n1125) );
  FD1S mem_reg_3__3_ ( .D(n610), .TI(mem_3__2_), .TE(test_se), .CP(n21), .Q(
        test_so3), .QN(n1124) );
  FD1S mem_reg_3__2_ ( .D(n609), .TI(mem_3__1_), .TE(test_se), .CP(n21), .Q(
        mem_3__2_), .QN(n1123) );
  FD1S mem_reg_3__1_ ( .D(n608), .TI(mem_3__0_), .TE(test_se), .CP(n21), .Q(
        mem_3__1_), .QN(n1122) );
  FD1S mem_reg_3__0_ ( .D(n643), .TI(mem_2__35_), .TE(test_se), .CP(n24), .Q(
        mem_3__0_), .QN(n1157) );
  FD1S mem_reg_2__35_ ( .D(n678), .TI(mem_2__34_), .TE(test_se), .CP(n18), .Q(
        mem_2__35_), .QN(n1192) );
  FD1S mem_reg_2__34_ ( .D(n677), .TI(mem_2__33_), .TE(test_se), .CP(n18), .Q(
        mem_2__34_), .QN(n1191) );
  FD1S mem_reg_2__33_ ( .D(n676), .TI(mem_2__32_), .TE(test_se), .CP(n17), .Q(
        mem_2__33_), .QN(n1190) );
  FD1S mem_reg_2__32_ ( .D(n675), .TI(mem_2__31_), .TE(test_se), .CP(n17), .Q(
        mem_2__32_), .QN(n1189) );
  FD1S mem_reg_2__31_ ( .D(n674), .TI(mem_2__30_), .TE(test_se), .CP(n17), .Q(
        mem_2__31_), .QN(n1188) );
  FD1S mem_reg_2__30_ ( .D(n673), .TI(mem_2__29_), .TE(test_se), .CP(n17), .Q(
        mem_2__30_), .QN(n1187) );
  FD1S mem_reg_2__29_ ( .D(n672), .TI(mem_2__28_), .TE(test_se), .CP(n17), .Q(
        mem_2__29_), .QN(n1186) );
  FD1S mem_reg_2__28_ ( .D(n671), .TI(mem_2__27_), .TE(test_se), .CP(n17), .Q(
        mem_2__28_), .QN(n1185) );
  FD1S mem_reg_2__27_ ( .D(n670), .TI(mem_2__26_), .TE(test_se), .CP(n17), .Q(
        mem_2__27_), .QN(n1184) );
  FD1S mem_reg_2__26_ ( .D(n669), .TI(mem_2__25_), .TE(test_se), .CP(n17), .Q(
        mem_2__26_), .QN(n1183) );
  FD1S mem_reg_2__25_ ( .D(n668), .TI(mem_2__24_), .TE(test_se), .CP(n17), .Q(
        mem_2__25_), .QN(n1182) );
  FD1S mem_reg_2__24_ ( .D(n667), .TI(mem_2__23_), .TE(test_se), .CP(n17), .Q(
        mem_2__24_), .QN(n1181) );
  FD1S mem_reg_2__23_ ( .D(n666), .TI(mem_2__22_), .TE(test_se), .CP(n17), .Q(
        mem_2__23_), .QN(n1180) );
  FD1S mem_reg_2__22_ ( .D(n665), .TI(mem_2__21_), .TE(test_se), .CP(n17), .Q(
        mem_2__22_), .QN(n1179) );
  FD1S mem_reg_2__21_ ( .D(n664), .TI(mem_2__20_), .TE(test_se), .CP(n16), .Q(
        mem_2__21_), .QN(n1178) );
  FD1S mem_reg_2__20_ ( .D(n663), .TI(mem_2__19_), .TE(test_se), .CP(n16), .Q(
        mem_2__20_), .QN(n1177) );
  FD1S mem_reg_2__19_ ( .D(n662), .TI(mem_2__18_), .TE(test_se), .CP(n16), .Q(
        mem_2__19_), .QN(n1176) );
  FD1S mem_reg_2__18_ ( .D(n661), .TI(mem_2__17_), .TE(test_se), .CP(n16), .Q(
        mem_2__18_), .QN(n1175) );
  FD1S mem_reg_2__17_ ( .D(n660), .TI(mem_2__16_), .TE(test_se), .CP(n16), .Q(
        mem_2__17_), .QN(n1174) );
  FD1S mem_reg_2__16_ ( .D(n659), .TI(mem_2__15_), .TE(test_se), .CP(n16), .Q(
        mem_2__16_), .QN(n1173) );
  FD1S mem_reg_2__15_ ( .D(n658), .TI(mem_2__14_), .TE(test_se), .CP(n16), .Q(
        mem_2__15_), .QN(n1172) );
  FD1S mem_reg_2__14_ ( .D(n657), .TI(mem_2__13_), .TE(test_se), .CP(n16), .Q(
        mem_2__14_), .QN(n1171) );
  FD1S mem_reg_2__13_ ( .D(n656), .TI(mem_2__12_), .TE(test_se), .CP(n16), .Q(
        mem_2__13_), .QN(n1170) );
  FD1S mem_reg_2__12_ ( .D(n655), .TI(mem_2__11_), .TE(test_se), .CP(n16), .Q(
        mem_2__12_), .QN(n1169) );
  FD1S mem_reg_2__11_ ( .D(n654), .TI(mem_2__10_), .TE(test_se), .CP(n16), .Q(
        mem_2__11_), .QN(n1168) );
  FD1S mem_reg_2__10_ ( .D(n653), .TI(mem_2__9_), .TE(test_se), .CP(n16), .Q(
        mem_2__10_), .QN(n1167) );
  FD1S mem_reg_2__9_ ( .D(n652), .TI(mem_2__8_), .TE(test_se), .CP(n15), .Q(
        mem_2__9_), .QN(n1166) );
  FD1S mem_reg_2__8_ ( .D(n651), .TI(mem_2__7_), .TE(test_se), .CP(n15), .Q(
        mem_2__8_), .QN(n1165) );
  FD1S mem_reg_2__7_ ( .D(n650), .TI(mem_2__6_), .TE(test_se), .CP(n15), .Q(
        mem_2__7_), .QN(n1164) );
  FD1S mem_reg_2__6_ ( .D(n649), .TI(mem_2__5_), .TE(test_se), .CP(n15), .Q(
        mem_2__6_), .QN(n1163) );
  FD1S mem_reg_2__5_ ( .D(n648), .TI(mem_2__4_), .TE(test_se), .CP(n15), .Q(
        mem_2__5_), .QN(n1162) );
  FD1S mem_reg_2__4_ ( .D(n647), .TI(mem_2__3_), .TE(test_se), .CP(n15), .Q(
        mem_2__4_), .QN(n1161) );
  FD1S mem_reg_2__3_ ( .D(n646), .TI(mem_2__2_), .TE(test_se), .CP(n15), .Q(
        mem_2__3_), .QN(n1160) );
  FD1S mem_reg_2__2_ ( .D(n645), .TI(mem_2__1_), .TE(test_se), .CP(n15), .Q(
        mem_2__2_), .QN(n1159) );
  FD1S mem_reg_2__1_ ( .D(n644), .TI(mem_2__0_), .TE(test_se), .CP(n15), .Q(
        mem_2__1_), .QN(n1158) );
  FD1S mem_reg_2__0_ ( .D(n679), .TI(mem_1__35_), .TE(test_se), .CP(n18), .Q(
        mem_2__0_), .QN(n1193) );
  FD1S mem_reg_1__35_ ( .D(n714), .TI(mem_1__34_), .TE(test_se), .CP(n21), .Q(
        mem_1__35_), .QN(n1228) );
  FD1S mem_reg_1__34_ ( .D(n713), .TI(mem_1__33_), .TE(test_se), .CP(n21), .Q(
        mem_1__34_), .QN(n1227) );
  FD1S mem_reg_1__33_ ( .D(n712), .TI(mem_1__32_), .TE(test_se), .CP(n20), .Q(
        mem_1__33_), .QN(n1226) );
  FD1S mem_reg_1__32_ ( .D(n711), .TI(mem_1__31_), .TE(test_se), .CP(n20), .Q(
        mem_1__32_), .QN(n1225) );
  FD1S mem_reg_1__31_ ( .D(n710), .TI(mem_1__30_), .TE(test_se), .CP(n20), .Q(
        mem_1__31_), .QN(n1224) );
  FD1S mem_reg_1__30_ ( .D(n709), .TI(mem_1__29_), .TE(test_se), .CP(n20), .Q(
        mem_1__30_), .QN(n1223) );
  FD1S mem_reg_1__29_ ( .D(n708), .TI(test_si3), .TE(test_se), .CP(n20), .Q(
        mem_1__29_), .QN(n1222) );
  FD1S mem_reg_1__28_ ( .D(n707), .TI(mem_1__27_), .TE(test_se), .CP(n20), .Q(
        test_so2), .QN(n1221) );
  FD1S mem_reg_1__27_ ( .D(n706), .TI(mem_1__26_), .TE(test_se), .CP(n20), .Q(
        mem_1__27_), .QN(n1220) );
  FD1S mem_reg_1__26_ ( .D(n705), .TI(mem_1__25_), .TE(test_se), .CP(n20), .Q(
        mem_1__26_), .QN(n1219) );
  FD1S mem_reg_1__25_ ( .D(n704), .TI(mem_1__24_), .TE(test_se), .CP(n20), .Q(
        mem_1__25_), .QN(n1218) );
  FD1S mem_reg_1__24_ ( .D(n703), .TI(mem_1__23_), .TE(test_se), .CP(n20), .Q(
        mem_1__24_), .QN(n1217) );
  FD1S mem_reg_1__23_ ( .D(n702), .TI(mem_1__22_), .TE(test_se), .CP(n20), .Q(
        mem_1__23_), .QN(n1216) );
  FD1S mem_reg_1__22_ ( .D(n701), .TI(mem_1__21_), .TE(test_se), .CP(n20), .Q(
        mem_1__22_), .QN(n1215) );
  FD1S mem_reg_1__21_ ( .D(n700), .TI(mem_1__20_), .TE(test_se), .CP(n19), .Q(
        mem_1__21_), .QN(n1214) );
  FD1S mem_reg_1__20_ ( .D(n699), .TI(mem_1__19_), .TE(test_se), .CP(n19), .Q(
        mem_1__20_), .QN(n1213) );
  FD1S mem_reg_1__19_ ( .D(n698), .TI(mem_1__18_), .TE(test_se), .CP(n19), .Q(
        mem_1__19_), .QN(n1212) );
  FD1S mem_reg_1__18_ ( .D(n697), .TI(mem_1__17_), .TE(test_se), .CP(n19), .Q(
        mem_1__18_), .QN(n1211) );
  FD1S mem_reg_1__17_ ( .D(n696), .TI(mem_1__16_), .TE(test_se), .CP(n19), .Q(
        mem_1__17_), .QN(n1210) );
  FD1S mem_reg_1__16_ ( .D(n695), .TI(mem_1__15_), .TE(test_se), .CP(n19), .Q(
        mem_1__16_), .QN(n1209) );
  FD1S mem_reg_1__15_ ( .D(n694), .TI(mem_1__14_), .TE(test_se), .CP(n19), .Q(
        mem_1__15_), .QN(n1208) );
  FD1S mem_reg_1__14_ ( .D(n693), .TI(mem_1__13_), .TE(test_se), .CP(n19), .Q(
        mem_1__14_), .QN(n1207) );
  FD1S mem_reg_1__13_ ( .D(n692), .TI(mem_1__12_), .TE(test_se), .CP(n19), .Q(
        mem_1__13_), .QN(n1206) );
  FD1S mem_reg_1__12_ ( .D(n691), .TI(mem_1__11_), .TE(test_se), .CP(n19), .Q(
        mem_1__12_), .QN(n1205) );
  FD1S mem_reg_1__11_ ( .D(n690), .TI(mem_1__10_), .TE(test_se), .CP(n19), .Q(
        mem_1__11_), .QN(n1204) );
  FD1S mem_reg_1__10_ ( .D(n689), .TI(mem_1__9_), .TE(test_se), .CP(n19), .Q(
        mem_1__10_), .QN(n1203) );
  FD1S mem_reg_1__9_ ( .D(n688), .TI(mem_1__8_), .TE(test_se), .CP(n18), .Q(
        mem_1__9_), .QN(n1202) );
  FD1S mem_reg_1__8_ ( .D(n687), .TI(mem_1__7_), .TE(test_se), .CP(n18), .Q(
        mem_1__8_), .QN(n1201) );
  FD1S mem_reg_1__7_ ( .D(n686), .TI(mem_1__6_), .TE(test_se), .CP(n18), .Q(
        mem_1__7_), .QN(n1200) );
  FD1S mem_reg_1__6_ ( .D(n685), .TI(mem_1__5_), .TE(test_se), .CP(n18), .Q(
        mem_1__6_), .QN(n1199) );
  FD1S mem_reg_1__5_ ( .D(n684), .TI(mem_1__4_), .TE(test_se), .CP(n18), .Q(
        mem_1__5_), .QN(n1198) );
  FD1S mem_reg_1__4_ ( .D(n683), .TI(mem_1__3_), .TE(test_se), .CP(n18), .Q(
        mem_1__4_), .QN(n1197) );
  FD1S mem_reg_1__3_ ( .D(n682), .TI(mem_1__2_), .TE(test_se), .CP(n18), .Q(
        mem_1__3_), .QN(n1196) );
  FD1S mem_reg_1__2_ ( .D(n681), .TI(mem_1__1_), .TE(test_se), .CP(n18), .Q(
        mem_1__2_), .QN(n1195) );
  FD1S mem_reg_1__1_ ( .D(n680), .TI(mem_1__0_), .TE(test_se), .CP(n18), .Q(
        mem_1__1_), .QN(n1194) );
  FD1S mem_reg_1__0_ ( .D(n715), .TI(mem_0__35_), .TE(test_se), .CP(n21), .Q(
        mem_1__0_), .QN(n1229) );
  FD1S mem_reg_0__35_ ( .D(n750), .TI(mem_0__34_), .TE(test_se), .CP(n30), .Q(
        mem_0__35_), .QN(n964) );
  FD1S mem_reg_0__34_ ( .D(n749), .TI(mem_0__33_), .TE(test_se), .CP(n30), .Q(
        mem_0__34_), .QN(n963) );
  FD1S mem_reg_0__33_ ( .D(n748), .TI(mem_0__32_), .TE(test_se), .CP(n30), .Q(
        mem_0__33_), .QN(n962) );
  FD1S mem_reg_0__32_ ( .D(n747), .TI(mem_0__31_), .TE(test_se), .CP(n30), .Q(
        mem_0__32_), .QN(n961) );
  FD1S mem_reg_0__31_ ( .D(n746), .TI(mem_0__30_), .TE(test_se), .CP(n29), .Q(
        mem_0__31_), .QN(n960) );
  FD1S mem_reg_0__30_ ( .D(n745), .TI(mem_0__29_), .TE(test_se), .CP(n29), .Q(
        mem_0__30_), .QN(n959) );
  FD1S mem_reg_0__29_ ( .D(n744), .TI(mem_0__28_), .TE(test_se), .CP(n29), .Q(
        mem_0__29_), .QN(n958) );
  FD1S mem_reg_0__28_ ( .D(n743), .TI(mem_0__27_), .TE(test_se), .CP(n29), .Q(
        mem_0__28_), .QN(n957) );
  FD1S mem_reg_0__27_ ( .D(n742), .TI(mem_0__26_), .TE(test_se), .CP(n29), .Q(
        mem_0__27_), .QN(n956) );
  FD1S mem_reg_0__26_ ( .D(n741), .TI(mem_0__25_), .TE(test_se), .CP(n29), .Q(
        mem_0__26_), .QN(n955) );
  FD1S mem_reg_0__25_ ( .D(n740), .TI(mem_0__24_), .TE(test_se), .CP(n29), .Q(
        mem_0__25_), .QN(n954) );
  FD1S mem_reg_0__24_ ( .D(n739), .TI(mem_0__23_), .TE(test_se), .CP(n29), .Q(
        mem_0__24_), .QN(n953) );
  FD1S mem_reg_0__23_ ( .D(n738), .TI(mem_0__22_), .TE(test_se), .CP(n29), .Q(
        mem_0__23_), .QN(n952) );
  FD1S mem_reg_0__22_ ( .D(n737), .TI(mem_0__21_), .TE(test_se), .CP(n29), .Q(
        mem_0__22_), .QN(n951) );
  FD1S mem_reg_0__21_ ( .D(n736), .TI(mem_0__20_), .TE(test_se), .CP(n29), .Q(
        mem_0__21_), .QN(n950) );
  FD1S mem_reg_0__20_ ( .D(n735), .TI(mem_0__19_), .TE(test_se), .CP(n29), .Q(
        mem_0__20_), .QN(n949) );
  FD1S mem_reg_0__19_ ( .D(n734), .TI(mem_0__18_), .TE(test_se), .CP(n28), .Q(
        mem_0__19_), .QN(n948) );
  FD1S mem_reg_0__18_ ( .D(n733), .TI(mem_0__17_), .TE(test_se), .CP(n28), .Q(
        mem_0__18_), .QN(n947) );
  FD1S mem_reg_0__17_ ( .D(n732), .TI(test_si2), .TE(test_se), .CP(n28), .Q(
        mem_0__17_), .QN(n946) );
  FD1S mem_reg_0__16_ ( .D(n731), .TI(mem_0__15_), .TE(test_se), .CP(n28), .Q(
        test_so1), .QN(n945) );
  FD1S mem_reg_0__15_ ( .D(n730), .TI(mem_0__14_), .TE(test_se), .CP(n28), .Q(
        mem_0__15_), .QN(n944) );
  FD1S mem_reg_0__14_ ( .D(n729), .TI(mem_0__13_), .TE(test_se), .CP(n28), .Q(
        mem_0__14_), .QN(n943) );
  FD1S mem_reg_0__13_ ( .D(n728), .TI(mem_0__12_), .TE(test_se), .CP(n28), .Q(
        mem_0__13_), .QN(n942) );
  FD1S mem_reg_0__12_ ( .D(n727), .TI(mem_0__11_), .TE(test_se), .CP(n28), .Q(
        mem_0__12_), .QN(n1241) );
  FD1S mem_reg_0__11_ ( .D(n726), .TI(mem_0__10_), .TE(test_se), .CP(n28), .Q(
        mem_0__11_), .QN(n1240) );
  FD1S mem_reg_0__10_ ( .D(n725), .TI(mem_0__9_), .TE(test_se), .CP(n28), .Q(
        mem_0__10_), .QN(n1239) );
  FD1S mem_reg_0__9_ ( .D(n724), .TI(mem_0__8_), .TE(test_se), .CP(n28), .Q(
        mem_0__9_), .QN(n1238) );
  FD1S mem_reg_0__8_ ( .D(n723), .TI(mem_0__7_), .TE(test_se), .CP(n28), .Q(
        mem_0__8_), .QN(n1237) );
  FD1S mem_reg_0__7_ ( .D(n722), .TI(mem_0__6_), .TE(test_se), .CP(n27), .Q(
        mem_0__7_), .QN(n1236) );
  FD1S mem_reg_0__6_ ( .D(n721), .TI(mem_0__5_), .TE(test_se), .CP(n27), .Q(
        mem_0__6_), .QN(n1235) );
  FD1S mem_reg_0__5_ ( .D(n720), .TI(mem_0__4_), .TE(test_se), .CP(n27), .Q(
        mem_0__5_), .QN(n1234) );
  FD1S mem_reg_0__4_ ( .D(n719), .TI(mem_0__3_), .TE(test_se), .CP(n27), .Q(
        mem_0__4_), .QN(n1233) );
  FD1S mem_reg_0__3_ ( .D(n718), .TI(mem_0__2_), .TE(test_se), .CP(n27), .Q(
        mem_0__3_), .QN(n1232) );
  FD1S mem_reg_0__2_ ( .D(n717), .TI(mem_0__1_), .TE(test_se), .CP(n27), .Q(
        mem_0__2_), .QN(n1231) );
  FD1S mem_reg_0__1_ ( .D(n716), .TI(mem_0__0_), .TE(test_se), .CP(n27), .Q(
        mem_0__1_), .QN(n1230) );
  FD1S mem_reg_0__0_ ( .D(n751), .TI(grey_wr_ptr[3]), .TE(test_se), .CP(n30), 
        .Q(mem_0__0_), .QN(n965) );
  FD2S grey_wr_ptr_reg_3_ ( .D(n461), .TI(grey_wr_ptr[2]), .TE(test_se), .CP(
        n12), .CD(wr_reset_n), .Q(grey_wr_ptr[3]), .QN(n976) );
  FD2S grey_wr_ptr_reg_2_ ( .D(n462), .TI(grey_wr_ptr[1]), .TE(test_se), .CP(
        n21), .CD(wr_reset_n), .Q(grey_wr_ptr[2]), .QN(n977) );
  FD2S grey_wr_ptr_reg_1_ ( .D(n459), .TI(grey_wr_ptr[0]), .TE(test_se), .CP(
        n21), .CD(wr_reset_n), .Q(grey_wr_ptr[1]), .QN(n974) );
  FD2S grey_wr_ptr_reg_0_ ( .D(n460), .TI(full), .TE(test_se), .CP(n5), .CD(
        wr_reset_n), .Q(grey_wr_ptr[0]), .QN(n975) );
  FD2S grey_rd_ptr_reg_1_ ( .D(n755), .TI(grey_rd_ptr_dly[0]), .TE(test_se), 
        .CP(rd_clk), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[1]), .QN(n966) );
  FD2S grey_rd_ptr_reg_3_ ( .D(n757), .TI(grey_rd_ptr_dly[2]), .TE(test_se), 
        .CP(rd_clk), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[3]), .QN(n967) );
  FD2S grey_rd_ptr_reg_2_ ( .D(n758), .TI(grey_rd_ptr_dly[1]), .TE(test_se), 
        .CP(rd_clk), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[2]), .QN(n968) );
  FD2S full_q_reg ( .D(n458), .TI(test_si1), .TE(test_se), .CP(n5), .CD(
        wr_reset_n), .Q(full), .QN(n972) );
  FD2S sync_rd_ptr_1_reg_0_ ( .D(sync_rd_ptr_0[0]), .TI(sync_rd_ptr_0[3]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[0]) );
  FD2S sync_rd_ptr_1_reg_2_ ( .D(sync_rd_ptr_0[2]), .TI(sync_rd_ptr_1[1]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[2]), .QN(n973) );
  FD2S sync_wr_ptr_1_reg_1_ ( .D(sync_wr_ptr_0[1]), .TI(sync_wr_ptr_1_0_), 
        .TE(test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(sync_wr_ptr_1_1_) );
  FD2S sync_wr_ptr_1_reg_0_ ( .D(sync_wr_ptr_0[0]), .TI(sync_wr_ptr_0[3]), 
        .TE(test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(sync_wr_ptr_1_0_) );
  FD2S wr_ptr_reg_0_ ( .D(n754), .TI(sync_rd_ptr_1[3]), .TE(test_se), .CP(n5), 
        .CD(wr_reset_n), .Q(n1242), .QN(n1) );
  FD2S wr_ptr_reg_3_ ( .D(n463), .TI(wr_ptr_2_), .TE(test_se), .CP(n12), .CD(
        wr_reset_n), .Q(test_so7) );
  FD2S grey_rd_ptr_reg_0_ ( .D(n756), .TI(test_si8), .TE(test_se), .CP(rd_clk), 
        .CD(rd_reset_n), .Q(grey_rd_ptr_dly[0]) );
  FD2S sync_rd_ptr_1_reg_1_ ( .D(sync_rd_ptr_0[1]), .TI(sync_rd_ptr_1[0]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[1]) );
  FD2S rd_ptr_reg_3_ ( .D(n759), .TI(N71), .TE(test_se), .CP(rd_clk), .CD(
        rd_reset_n), .Q(rd_ptr_3_1), .QN(n4) );
  FD2S sync_wr_ptr_1_reg_3_ ( .D(sync_wr_ptr_0[3]), .TI(n1244), .TE(test_se), 
        .CP(rd_clk), .CD(rd_reset_n), .Q(test_so8) );
  FD2S rd_ptr_reg_1_ ( .D(n761), .TI(N69), .TE(test_se), .CP(rd_clk), .CD(
        rd_reset_n), .Q(N70), .QN(n969) );
  FD2S rd_ptr_reg_2_ ( .D(n760), .TI(N70), .TE(test_se), .CP(rd_clk), .CD(
        rd_reset_n), .Q(N71), .QN(n360) );
  FD2S sync_rd_ptr_1_reg_3_ ( .D(sync_rd_ptr_0[3]), .TI(sync_rd_ptr_1[2]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_1[3]) );
  FD2S rd_ptr_reg_0_ ( .D(n762), .TI(grey_rd_ptr_dly[3]), .TE(test_se), .CP(
        rd_clk), .CD(rd_reset_n), .Q(N69), .QN(n970) );
  FD2S wr_ptr_reg_1_ ( .D(n753), .TI(n1242), .TE(test_se), .CP(n5), .CD(
        wr_reset_n), .Q(wr_ptr_1_), .QN(n3) );
  FD2S wr_ptr_reg_2_ ( .D(n752), .TI(wr_ptr_1_), .TE(test_se), .CP(n6), .CD(
        wr_reset_n), .Q(wr_ptr_2_), .QN(n2) );
  FD2S sync_rd_ptr_0_reg_0_ ( .D(grey_rd_ptr_dly[0]), .TI(mem_7__35_), .TE(
        test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[0]) );
  FD2S sync_rd_ptr_0_reg_1_ ( .D(grey_rd_ptr_dly[1]), .TI(sync_rd_ptr_0[0]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[1]) );
  FD2S sync_rd_ptr_0_reg_3_ ( .D(grey_rd_ptr_dly[3]), .TI(sync_rd_ptr_0[2]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[3]) );
  FD2S sync_rd_ptr_0_reg_2_ ( .D(grey_rd_ptr_dly[2]), .TI(sync_rd_ptr_0[1]), 
        .TE(test_se), .CP(n5), .CD(wr_reset_n), .Q(sync_rd_ptr_0[2]) );
  FD2S sync_wr_ptr_0_reg_3_ ( .D(grey_wr_ptr[3]), .TI(sync_wr_ptr_0[2]), .TE(
        test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(sync_wr_ptr_0[3]) );
  FD2S sync_wr_ptr_0_reg_2_ ( .D(grey_wr_ptr[2]), .TI(sync_wr_ptr_0[1]), .TE(
        test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(sync_wr_ptr_0[2]) );
  FD2S sync_wr_ptr_0_reg_1_ ( .D(grey_wr_ptr[1]), .TI(sync_wr_ptr_0[0]), .TE(
        test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(sync_wr_ptr_0[1]) );
  FD2S sync_wr_ptr_0_reg_0_ ( .D(grey_wr_ptr[0]), .TI(rd_ptr_3_1), .TE(test_se), .CP(rd_clk), .CD(rd_reset_n), .Q(sync_wr_ptr_0[0]) );
  IVP U324 ( .A(n31), .Z(n28) );
  IVP U325 ( .A(n31), .Z(n29) );
  IVP U326 ( .A(n34), .Z(n19) );
  IVP U327 ( .A(n34), .Z(n20) );
  IVP U328 ( .A(n356), .Z(n16) );
  IVP U329 ( .A(n356), .Z(n17) );
  IVP U330 ( .A(n356), .Z(n18) );
  IVP U331 ( .A(n33), .Z(n22) );
  IVP U332 ( .A(n33), .Z(n23) );
  IVP U333 ( .A(n33), .Z(n24) );
  IVP U334 ( .A(n32), .Z(n25) );
  IVP U335 ( .A(n32), .Z(n26) );
  IVP U336 ( .A(n32), .Z(n27) );
  IVP U337 ( .A(n359), .Z(n7) );
  IVP U338 ( .A(n359), .Z(n8) );
  IVP U339 ( .A(n359), .Z(n9) );
  IVP U340 ( .A(n358), .Z(n10) );
  IVP U341 ( .A(n358), .Z(n11) );
  IVP U342 ( .A(n357), .Z(n13) );
  IVP U343 ( .A(n357), .Z(n14) );
  IVP U344 ( .A(n357), .Z(n15) );
  IVP U345 ( .A(n34), .Z(n21) );
  IVP U346 ( .A(n358), .Z(n12) );
  IVP U347 ( .A(n361), .Z(n6) );
  IVP U348 ( .A(n361), .Z(n5) );
  IVP U349 ( .A(n31), .Z(n30) );
  IVP U350 ( .A(n364), .Z(n31) );
  IVP U351 ( .A(n363), .Z(n356) );
  IVP U352 ( .A(n364), .Z(n33) );
  IVP U353 ( .A(n364), .Z(n32) );
  IVP U354 ( .A(n362), .Z(n359) );
  IVP U355 ( .A(n363), .Z(n357) );
  IVP U356 ( .A(n363), .Z(n34) );
  IVP U357 ( .A(n362), .Z(n358) );
  IVP U358 ( .A(n362), .Z(n361) );
  IVP U359 ( .A(n365), .Z(n364) );
  IVP U360 ( .A(n365), .Z(n363) );
  IVP U361 ( .A(n365), .Z(n362) );
  IVP U362 ( .A(wr_clk), .Z(n365) );
  ND2 U363 ( .A(N71), .B(n969), .Z(n366) );
  NR2 U364 ( .A(n366), .B(n970), .Z(n816) );
  ND2 U365 ( .A(N71), .B(N70), .Z(n367) );
  NR2 U366 ( .A(n970), .B(n367), .Z(n815) );
  AO2 U367 ( .A(mem_5__0_), .B(n816), .C(test_so6), .D(n815), .Z(n373) );
  ND2 U368 ( .A(n969), .B(n360), .Z(n368) );
  NR2 U369 ( .A(n368), .B(n970), .Z(n818) );
  ND2 U370 ( .A(N70), .B(n360), .Z(n369) );
  NR2 U371 ( .A(n369), .B(n970), .Z(n817) );
  AO2 U372 ( .A(mem_1__0_), .B(n818), .C(mem_3__0_), .D(n817), .Z(n372) );
  NR2 U373 ( .A(n366), .B(N69), .Z(n820) );
  NR2 U374 ( .A(n367), .B(N69), .Z(n819) );
  AO2 U375 ( .A(mem_4__0_), .B(n820), .C(mem_6__0_), .D(n819), .Z(n371) );
  NR2 U376 ( .A(n368), .B(N69), .Z(n822) );
  NR2 U377 ( .A(n369), .B(N69), .Z(n821) );
  AO2 U378 ( .A(mem_0__0_), .B(n822), .C(mem_2__0_), .D(n821), .Z(n370) );
  ND4 U379 ( .A(n373), .B(n372), .C(n371), .D(n370), .Z(rd_data[0]) );
  AO2 U380 ( .A(mem_5__1_), .B(n816), .C(mem_7__1_), .D(n815), .Z(n377) );
  AO2 U381 ( .A(mem_1__1_), .B(n818), .C(mem_3__1_), .D(n817), .Z(n376) );
  AO2 U382 ( .A(mem_4__1_), .B(n820), .C(mem_6__1_), .D(n819), .Z(n375) );
  AO2 U383 ( .A(mem_0__1_), .B(n822), .C(mem_2__1_), .D(n821), .Z(n374) );
  ND4 U384 ( .A(n377), .B(n376), .C(n375), .D(n374), .Z(rd_data[1]) );
  AO2 U385 ( .A(mem_5__2_), .B(n816), .C(mem_7__2_), .D(n815), .Z(n381) );
  AO2 U386 ( .A(mem_1__2_), .B(n818), .C(mem_3__2_), .D(n817), .Z(n380) );
  AO2 U387 ( .A(mem_4__2_), .B(n820), .C(mem_6__2_), .D(n819), .Z(n379) );
  AO2 U388 ( .A(mem_0__2_), .B(n822), .C(mem_2__2_), .D(n821), .Z(n378) );
  ND4 U389 ( .A(n381), .B(n380), .C(n379), .D(n378), .Z(rd_data[2]) );
  AO2 U390 ( .A(mem_5__3_), .B(n816), .C(mem_7__3_), .D(n815), .Z(n385) );
  AO2 U391 ( .A(mem_1__3_), .B(n818), .C(test_so3), .D(n817), .Z(n384) );
  AO2 U392 ( .A(mem_4__3_), .B(n820), .C(mem_6__3_), .D(n819), .Z(n383) );
  AO2 U393 ( .A(mem_0__3_), .B(n822), .C(mem_2__3_), .D(n821), .Z(n382) );
  ND4 U394 ( .A(n385), .B(n384), .C(n383), .D(n382), .Z(rd_data[3]) );
  AO2 U395 ( .A(mem_5__4_), .B(n816), .C(mem_7__4_), .D(n815), .Z(n389) );
  AO2 U396 ( .A(mem_1__4_), .B(n818), .C(mem_3__4_), .D(n817), .Z(n388) );
  AO2 U397 ( .A(mem_4__4_), .B(n820), .C(mem_6__4_), .D(n819), .Z(n387) );
  AO2 U398 ( .A(mem_0__4_), .B(n822), .C(mem_2__4_), .D(n821), .Z(n386) );
  ND4 U399 ( .A(n389), .B(n388), .C(n387), .D(n386), .Z(rd_data[4]) );
  AO2 U400 ( .A(mem_5__5_), .B(n816), .C(mem_7__5_), .D(n815), .Z(n393) );
  AO2 U401 ( .A(mem_1__5_), .B(n818), .C(mem_3__5_), .D(n817), .Z(n392) );
  AO2 U402 ( .A(mem_4__5_), .B(n820), .C(mem_6__5_), .D(n819), .Z(n391) );
  AO2 U403 ( .A(mem_0__5_), .B(n822), .C(mem_2__5_), .D(n821), .Z(n390) );
  ND4 U404 ( .A(n393), .B(n392), .C(n391), .D(n390), .Z(rd_data[5]) );
  AO2 U405 ( .A(mem_5__6_), .B(n816), .C(mem_7__6_), .D(n815), .Z(n397) );
  AO2 U406 ( .A(mem_1__6_), .B(n818), .C(mem_3__6_), .D(n817), .Z(n396) );
  AO2 U407 ( .A(mem_4__6_), .B(n820), .C(mem_6__6_), .D(n819), .Z(n395) );
  AO2 U408 ( .A(mem_0__6_), .B(n822), .C(mem_2__6_), .D(n821), .Z(n394) );
  ND4 U409 ( .A(n397), .B(n396), .C(n395), .D(n394), .Z(rd_data[6]) );
  AO2 U410 ( .A(mem_5__7_), .B(n816), .C(mem_7__7_), .D(n815), .Z(n401) );
  AO2 U411 ( .A(mem_1__7_), .B(n818), .C(mem_3__7_), .D(n817), .Z(n400) );
  AO2 U412 ( .A(mem_4__7_), .B(n820), .C(mem_6__7_), .D(n819), .Z(n399) );
  AO2 U413 ( .A(mem_0__7_), .B(n822), .C(mem_2__7_), .D(n821), .Z(n398) );
  ND4 U414 ( .A(n401), .B(n400), .C(n399), .D(n398), .Z(rd_data[7]) );
  AO2 U415 ( .A(mem_5__8_), .B(n816), .C(mem_7__8_), .D(n815), .Z(n405) );
  AO2 U416 ( .A(mem_1__8_), .B(n818), .C(mem_3__8_), .D(n817), .Z(n404) );
  AO2 U417 ( .A(mem_4__8_), .B(n820), .C(mem_6__8_), .D(n819), .Z(n403) );
  AO2 U418 ( .A(mem_0__8_), .B(n822), .C(mem_2__8_), .D(n821), .Z(n402) );
  ND4 U419 ( .A(n405), .B(n404), .C(n403), .D(n402), .Z(rd_data[8]) );
  AO2 U420 ( .A(mem_5__9_), .B(n816), .C(mem_7__9_), .D(n815), .Z(n409) );
  AO2 U421 ( .A(mem_1__9_), .B(n818), .C(mem_3__9_), .D(n817), .Z(n408) );
  AO2 U422 ( .A(mem_4__9_), .B(n820), .C(mem_6__9_), .D(n819), .Z(n407) );
  AO2 U423 ( .A(mem_0__9_), .B(n822), .C(mem_2__9_), .D(n821), .Z(n406) );
  ND4 U424 ( .A(n409), .B(n408), .C(n407), .D(n406), .Z(rd_data[9]) );
  AO2 U425 ( .A(mem_5__10_), .B(n816), .C(mem_7__10_), .D(n815), .Z(n413) );
  AO2 U426 ( .A(mem_1__10_), .B(n818), .C(mem_3__10_), .D(n817), .Z(n412) );
  AO2 U427 ( .A(mem_4__10_), .B(n820), .C(mem_6__10_), .D(n819), .Z(n411) );
  AO2 U428 ( .A(mem_0__10_), .B(n822), .C(mem_2__10_), .D(n821), .Z(n410) );
  ND4 U429 ( .A(n413), .B(n412), .C(n411), .D(n410), .Z(rd_data[10]) );
  AO2 U430 ( .A(mem_5__11_), .B(n816), .C(mem_7__11_), .D(n815), .Z(n417) );
  AO2 U431 ( .A(mem_1__11_), .B(n818), .C(mem_3__11_), .D(n817), .Z(n416) );
  AO2 U432 ( .A(mem_4__11_), .B(n820), .C(mem_6__11_), .D(n819), .Z(n415) );
  AO2 U433 ( .A(mem_0__11_), .B(n822), .C(mem_2__11_), .D(n821), .Z(n414) );
  ND4 U434 ( .A(n417), .B(n416), .C(n415), .D(n414), .Z(rd_data[11]) );
  AO2 U435 ( .A(mem_5__12_), .B(n816), .C(mem_7__12_), .D(n815), .Z(n421) );
  AO2 U436 ( .A(mem_1__12_), .B(n818), .C(mem_3__12_), .D(n817), .Z(n420) );
  AO2 U437 ( .A(mem_4__12_), .B(n820), .C(mem_6__12_), .D(n819), .Z(n419) );
  AO2 U438 ( .A(mem_0__12_), .B(n822), .C(mem_2__12_), .D(n821), .Z(n418) );
  ND4 U439 ( .A(n421), .B(n420), .C(n419), .D(n418), .Z(rd_data[12]) );
  AO2 U440 ( .A(mem_5__13_), .B(n816), .C(mem_7__13_), .D(n815), .Z(n425) );
  AO2 U441 ( .A(mem_1__13_), .B(n818), .C(mem_3__13_), .D(n817), .Z(n424) );
  AO2 U442 ( .A(mem_4__13_), .B(n820), .C(mem_6__13_), .D(n819), .Z(n423) );
  AO2 U443 ( .A(mem_0__13_), .B(n822), .C(mem_2__13_), .D(n821), .Z(n422) );
  ND4 U444 ( .A(n425), .B(n424), .C(n423), .D(n422), .Z(rd_data[13]) );
  AO2 U445 ( .A(mem_5__14_), .B(n816), .C(mem_7__14_), .D(n815), .Z(n429) );
  AO2 U446 ( .A(mem_1__14_), .B(n818), .C(mem_3__14_), .D(n817), .Z(n428) );
  AO2 U447 ( .A(test_so4), .B(n820), .C(mem_6__14_), .D(n819), .Z(n427) );
  AO2 U448 ( .A(mem_0__14_), .B(n822), .C(mem_2__14_), .D(n821), .Z(n426) );
  ND4 U449 ( .A(n429), .B(n428), .C(n427), .D(n426), .Z(rd_data[14]) );
  AO2 U450 ( .A(mem_5__15_), .B(n816), .C(mem_7__15_), .D(n815), .Z(n433) );
  AO2 U451 ( .A(mem_1__15_), .B(n818), .C(mem_3__15_), .D(n817), .Z(n432) );
  AO2 U452 ( .A(mem_4__15_), .B(n820), .C(mem_6__15_), .D(n819), .Z(n431) );
  AO2 U453 ( .A(mem_0__15_), .B(n822), .C(mem_2__15_), .D(n821), .Z(n430) );
  ND4 U454 ( .A(n433), .B(n432), .C(n431), .D(n430), .Z(rd_data[15]) );
  AO2 U455 ( .A(mem_5__16_), .B(n816), .C(mem_7__16_), .D(n815), .Z(n437) );
  AO2 U456 ( .A(mem_1__16_), .B(n818), .C(mem_3__16_), .D(n817), .Z(n436) );
  AO2 U457 ( .A(mem_4__16_), .B(n820), .C(mem_6__16_), .D(n819), .Z(n435) );
  AO2 U458 ( .A(test_so1), .B(n822), .C(mem_2__16_), .D(n821), .Z(n434) );
  ND4 U459 ( .A(n437), .B(n436), .C(n435), .D(n434), .Z(rd_data[16]) );
  AO2 U460 ( .A(mem_5__17_), .B(n816), .C(mem_7__17_), .D(n815), .Z(n441) );
  AO2 U461 ( .A(mem_1__17_), .B(n818), .C(mem_3__17_), .D(n817), .Z(n440) );
  AO2 U462 ( .A(mem_4__17_), .B(n820), .C(mem_6__17_), .D(n819), .Z(n439) );
  AO2 U463 ( .A(mem_0__17_), .B(n822), .C(mem_2__17_), .D(n821), .Z(n438) );
  ND4 U464 ( .A(n441), .B(n440), .C(n439), .D(n438), .Z(rd_data[17]) );
  AO2 U465 ( .A(mem_5__18_), .B(n816), .C(mem_7__18_), .D(n815), .Z(n445) );
  AO2 U466 ( .A(mem_1__18_), .B(n818), .C(mem_3__18_), .D(n817), .Z(n444) );
  AO2 U467 ( .A(mem_4__18_), .B(n820), .C(mem_6__18_), .D(n819), .Z(n443) );
  AO2 U468 ( .A(mem_0__18_), .B(n822), .C(mem_2__18_), .D(n821), .Z(n442) );
  ND4 U469 ( .A(n445), .B(n444), .C(n443), .D(n442), .Z(rd_data[18]) );
  AO2 U470 ( .A(mem_5__19_), .B(n816), .C(mem_7__19_), .D(n815), .Z(n449) );
  AO2 U471 ( .A(mem_1__19_), .B(n818), .C(mem_3__19_), .D(n817), .Z(n448) );
  AO2 U472 ( .A(mem_4__19_), .B(n820), .C(mem_6__19_), .D(n819), .Z(n447) );
  AO2 U473 ( .A(mem_0__19_), .B(n822), .C(mem_2__19_), .D(n821), .Z(n446) );
  ND4 U474 ( .A(n449), .B(n448), .C(n447), .D(n446), .Z(rd_data[19]) );
  AO2 U475 ( .A(mem_5__20_), .B(n816), .C(mem_7__20_), .D(n815), .Z(n453) );
  AO2 U476 ( .A(mem_1__20_), .B(n818), .C(mem_3__20_), .D(n817), .Z(n452) );
  AO2 U477 ( .A(mem_4__20_), .B(n820), .C(mem_6__20_), .D(n819), .Z(n451) );
  AO2 U478 ( .A(mem_0__20_), .B(n822), .C(mem_2__20_), .D(n821), .Z(n450) );
  ND4 U479 ( .A(n453), .B(n452), .C(n451), .D(n450), .Z(rd_data[20]) );
  AO2 U480 ( .A(mem_5__21_), .B(n816), .C(mem_7__21_), .D(n815), .Z(n457) );
  AO2 U481 ( .A(mem_1__21_), .B(n818), .C(mem_3__21_), .D(n817), .Z(n456) );
  AO2 U482 ( .A(mem_4__21_), .B(n820), .C(mem_6__21_), .D(n819), .Z(n455) );
  AO2 U483 ( .A(mem_0__21_), .B(n822), .C(mem_2__21_), .D(n821), .Z(n454) );
  ND4 U484 ( .A(n457), .B(n456), .C(n455), .D(n454), .Z(rd_data[21]) );
  AO2 U485 ( .A(mem_5__22_), .B(n816), .C(mem_7__22_), .D(n815), .Z(n766) );
  AO2 U486 ( .A(mem_1__22_), .B(n818), .C(mem_3__22_), .D(n817), .Z(n765) );
  AO2 U487 ( .A(mem_4__22_), .B(n820), .C(mem_6__22_), .D(n819), .Z(n764) );
  AO2 U488 ( .A(mem_0__22_), .B(n822), .C(mem_2__22_), .D(n821), .Z(n763) );
  ND4 U489 ( .A(n766), .B(n765), .C(n764), .D(n763), .Z(rd_data[22]) );
  AO2 U490 ( .A(mem_5__23_), .B(n816), .C(mem_7__23_), .D(n815), .Z(n770) );
  AO2 U491 ( .A(mem_1__23_), .B(n818), .C(mem_3__23_), .D(n817), .Z(n769) );
  AO2 U492 ( .A(mem_4__23_), .B(n820), .C(mem_6__23_), .D(n819), .Z(n768) );
  AO2 U493 ( .A(mem_0__23_), .B(n822), .C(mem_2__23_), .D(n821), .Z(n767) );
  ND4 U494 ( .A(n770), .B(n769), .C(n768), .D(n767), .Z(rd_data[23]) );
  AO2 U495 ( .A(mem_5__24_), .B(n816), .C(mem_7__24_), .D(n815), .Z(n774) );
  AO2 U496 ( .A(mem_1__24_), .B(n818), .C(mem_3__24_), .D(n817), .Z(n773) );
  AO2 U497 ( .A(mem_4__24_), .B(n820), .C(mem_6__24_), .D(n819), .Z(n772) );
  AO2 U498 ( .A(mem_0__24_), .B(n822), .C(mem_2__24_), .D(n821), .Z(n771) );
  ND4 U499 ( .A(n774), .B(n773), .C(n772), .D(n771), .Z(rd_data[24]) );
  AO2 U500 ( .A(test_so5), .B(n816), .C(mem_7__25_), .D(n815), .Z(n778) );
  AO2 U501 ( .A(mem_1__25_), .B(n818), .C(mem_3__25_), .D(n817), .Z(n777) );
  AO2 U502 ( .A(mem_4__25_), .B(n820), .C(mem_6__25_), .D(n819), .Z(n776) );
  AO2 U503 ( .A(mem_0__25_), .B(n822), .C(mem_2__25_), .D(n821), .Z(n775) );
  ND4 U504 ( .A(n778), .B(n777), .C(n776), .D(n775), .Z(rd_data[25]) );
  AO2 U505 ( .A(mem_5__26_), .B(n816), .C(mem_7__26_), .D(n815), .Z(n782) );
  AO2 U506 ( .A(mem_1__26_), .B(n818), .C(mem_3__26_), .D(n817), .Z(n781) );
  AO2 U507 ( .A(mem_4__26_), .B(n820), .C(mem_6__26_), .D(n819), .Z(n780) );
  AO2 U508 ( .A(mem_0__26_), .B(n822), .C(mem_2__26_), .D(n821), .Z(n779) );
  ND4 U509 ( .A(n782), .B(n781), .C(n780), .D(n779), .Z(rd_data[26]) );
  AO2 U510 ( .A(mem_5__27_), .B(n816), .C(mem_7__27_), .D(n815), .Z(n786) );
  AO2 U511 ( .A(mem_1__27_), .B(n818), .C(mem_3__27_), .D(n817), .Z(n785) );
  AO2 U512 ( .A(mem_4__27_), .B(n820), .C(mem_6__27_), .D(n819), .Z(n784) );
  AO2 U513 ( .A(mem_0__27_), .B(n822), .C(mem_2__27_), .D(n821), .Z(n783) );
  ND4 U514 ( .A(n786), .B(n785), .C(n784), .D(n783), .Z(rd_data[27]) );
  AO2 U515 ( .A(mem_5__28_), .B(n816), .C(mem_7__28_), .D(n815), .Z(n790) );
  AO2 U516 ( .A(test_so2), .B(n818), .C(mem_3__28_), .D(n817), .Z(n789) );
  AO2 U517 ( .A(mem_4__28_), .B(n820), .C(mem_6__28_), .D(n819), .Z(n788) );
  AO2 U518 ( .A(mem_0__28_), .B(n822), .C(mem_2__28_), .D(n821), .Z(n787) );
  ND4 U519 ( .A(n790), .B(n789), .C(n788), .D(n787), .Z(rd_data[28]) );
  AO2 U520 ( .A(mem_5__29_), .B(n816), .C(mem_7__29_), .D(n815), .Z(n794) );
  AO2 U521 ( .A(mem_1__29_), .B(n818), .C(mem_3__29_), .D(n817), .Z(n793) );
  AO2 U522 ( .A(mem_4__29_), .B(n820), .C(mem_6__29_), .D(n819), .Z(n792) );
  AO2 U523 ( .A(mem_0__29_), .B(n822), .C(mem_2__29_), .D(n821), .Z(n791) );
  ND4 U524 ( .A(n794), .B(n793), .C(n792), .D(n791), .Z(rd_data[29]) );
  AO2 U525 ( .A(mem_5__30_), .B(n816), .C(mem_7__30_), .D(n815), .Z(n798) );
  AO2 U526 ( .A(mem_1__30_), .B(n818), .C(mem_3__30_), .D(n817), .Z(n797) );
  AO2 U527 ( .A(mem_4__30_), .B(n820), .C(mem_6__30_), .D(n819), .Z(n796) );
  AO2 U528 ( .A(mem_0__30_), .B(n822), .C(mem_2__30_), .D(n821), .Z(n795) );
  ND4 U529 ( .A(n798), .B(n797), .C(n796), .D(n795), .Z(rd_data[30]) );
  AO2 U530 ( .A(mem_5__31_), .B(n816), .C(mem_7__31_), .D(n815), .Z(n802) );
  AO2 U531 ( .A(mem_1__31_), .B(n818), .C(mem_3__31_), .D(n817), .Z(n801) );
  AO2 U532 ( .A(mem_4__31_), .B(n820), .C(mem_6__31_), .D(n819), .Z(n800) );
  AO2 U533 ( .A(mem_0__31_), .B(n822), .C(mem_2__31_), .D(n821), .Z(n799) );
  ND4 U534 ( .A(n802), .B(n801), .C(n800), .D(n799), .Z(rd_data[31]) );
  AO2 U535 ( .A(mem_5__32_), .B(n816), .C(mem_7__32_), .D(n815), .Z(n806) );
  AO2 U536 ( .A(mem_1__32_), .B(n818), .C(mem_3__32_), .D(n817), .Z(n805) );
  AO2 U537 ( .A(mem_4__32_), .B(n820), .C(mem_6__32_), .D(n819), .Z(n804) );
  AO2 U538 ( .A(mem_0__32_), .B(n822), .C(mem_2__32_), .D(n821), .Z(n803) );
  ND4 U539 ( .A(n806), .B(n805), .C(n804), .D(n803), .Z(rd_data[32]) );
  AO2 U540 ( .A(mem_5__33_), .B(n816), .C(mem_7__33_), .D(n815), .Z(n810) );
  AO2 U541 ( .A(mem_1__33_), .B(n818), .C(mem_3__33_), .D(n817), .Z(n809) );
  AO2 U542 ( .A(mem_4__33_), .B(n820), .C(mem_6__33_), .D(n819), .Z(n808) );
  AO2 U543 ( .A(mem_0__33_), .B(n822), .C(mem_2__33_), .D(n821), .Z(n807) );
  ND4 U544 ( .A(n810), .B(n809), .C(n808), .D(n807), .Z(rd_data[33]) );
  AO2 U545 ( .A(mem_5__34_), .B(n816), .C(mem_7__34_), .D(n815), .Z(n814) );
  AO2 U546 ( .A(mem_1__34_), .B(n818), .C(mem_3__34_), .D(n817), .Z(n813) );
  AO2 U547 ( .A(mem_4__34_), .B(n820), .C(mem_6__34_), .D(n819), .Z(n812) );
  AO2 U548 ( .A(mem_0__34_), .B(n822), .C(mem_2__34_), .D(n821), .Z(n811) );
  ND4 U549 ( .A(n814), .B(n813), .C(n812), .D(n811), .Z(rd_data[34]) );
  AO2 U550 ( .A(mem_5__35_), .B(n816), .C(mem_7__35_), .D(n815), .Z(n826) );
  AO2 U551 ( .A(mem_1__35_), .B(n818), .C(mem_3__35_), .D(n817), .Z(n825) );
  AO2 U552 ( .A(mem_4__35_), .B(n820), .C(mem_6__35_), .D(n819), .Z(n824) );
  AO2 U553 ( .A(mem_0__35_), .B(n822), .C(mem_2__35_), .D(n821), .Z(n823) );
  ND4 U554 ( .A(n826), .B(n825), .C(n824), .D(n823), .Z(rd_data[35]) );
  EN U555 ( .A(n970), .B(rd_en), .Z(n762) );
  AO7 U556 ( .A(rd_en), .B(n969), .C(n827), .Z(n761) );
  IV U557 ( .A(n828), .Z(n760) );
  AO6 U558 ( .A(n829), .B(N71), .C(n830), .Z(n828) );
  AO7 U559 ( .A(rd_en), .B(n4), .C(n831), .Z(n759) );
  AO7 U560 ( .A(rd_en), .B(n968), .C(n832), .Z(n758) );
  AO2 U561 ( .A(n833), .B(n834), .C(n830), .D(n835), .Z(n832) );
  AO7 U562 ( .A(rd_en), .B(n967), .C(n831), .Z(n757) );
  IV U563 ( .A(n833), .Z(n831) );
  NR2 U564 ( .A(n829), .B(n835), .Z(n833) );
  EO U565 ( .A(n836), .B(rd_ptr_3_1), .Z(n835) );
  ND2 U566 ( .A(n837), .B(N71), .Z(n836) );
  AO7 U567 ( .A(n970), .B(n827), .C(n838), .Z(n756) );
  MUX21L U568 ( .A(n839), .B(grey_rd_ptr_dly[0]), .S(n829), .Z(n838) );
  NR2 U569 ( .A(n840), .B(N69), .Z(n839) );
  AO7 U570 ( .A(rd_en), .B(n966), .C(n841), .Z(n755) );
  AO2 U571 ( .A(n842), .B(n834), .C(n830), .D(n843), .Z(n841) );
  IV U572 ( .A(n840), .Z(n843) );
  NR2 U573 ( .A(n834), .B(n829), .Z(n830) );
  IV U574 ( .A(rd_en), .Z(n829) );
  EO U575 ( .A(n360), .B(n837), .Z(n834) );
  IV U576 ( .A(n827), .Z(n842) );
  ND2 U577 ( .A(n840), .B(rd_en), .Z(n827) );
  AO6 U578 ( .A(n970), .B(n969), .C(n837), .Z(n840) );
  AO7 U579 ( .A(wr_en), .B(n1), .C(n844), .Z(n754) );
  IV U580 ( .A(n845), .Z(n844) );
  IV U581 ( .A(n846), .Z(n753) );
  AO6 U582 ( .A(n847), .B(wr_ptr_1_), .C(n848), .Z(n846) );
  IV U583 ( .A(n849), .Z(n752) );
  AO6 U584 ( .A(n847), .B(wr_ptr_2_), .C(n850), .Z(n849) );
  MUX21L U585 ( .A(n965), .B(n851), .S(n852), .Z(n751) );
  MUX21L U586 ( .A(n964), .B(n853), .S(n852), .Z(n750) );
  MUX21L U587 ( .A(n963), .B(n854), .S(n852), .Z(n749) );
  MUX21L U588 ( .A(n962), .B(n855), .S(n852), .Z(n748) );
  MUX21L U589 ( .A(n961), .B(n856), .S(n852), .Z(n747) );
  MUX21L U590 ( .A(n960), .B(n857), .S(n852), .Z(n746) );
  MUX21L U591 ( .A(n959), .B(n858), .S(n852), .Z(n745) );
  MUX21L U592 ( .A(n958), .B(n859), .S(n852), .Z(n744) );
  MUX21L U593 ( .A(n957), .B(n860), .S(n852), .Z(n743) );
  MUX21L U594 ( .A(n956), .B(n861), .S(n852), .Z(n742) );
  MUX21L U595 ( .A(n955), .B(n862), .S(n852), .Z(n741) );
  MUX21L U596 ( .A(n954), .B(n863), .S(n852), .Z(n740) );
  MUX21L U597 ( .A(n953), .B(n864), .S(n852), .Z(n739) );
  MUX21L U598 ( .A(n952), .B(n865), .S(n852), .Z(n738) );
  MUX21L U599 ( .A(n951), .B(n866), .S(n852), .Z(n737) );
  MUX21L U600 ( .A(n950), .B(n867), .S(n852), .Z(n736) );
  MUX21L U601 ( .A(n949), .B(n868), .S(n852), .Z(n735) );
  MUX21L U602 ( .A(n948), .B(n869), .S(n852), .Z(n734) );
  MUX21L U603 ( .A(n947), .B(n870), .S(n852), .Z(n733) );
  MUX21L U604 ( .A(n946), .B(n871), .S(n852), .Z(n732) );
  MUX21L U605 ( .A(n945), .B(n872), .S(n852), .Z(n731) );
  MUX21L U606 ( .A(n944), .B(n873), .S(n852), .Z(n730) );
  MUX21L U607 ( .A(n943), .B(n874), .S(n852), .Z(n729) );
  MUX21L U608 ( .A(n942), .B(n875), .S(n852), .Z(n728) );
  MUX21L U609 ( .A(n1241), .B(n876), .S(n852), .Z(n727) );
  MUX21L U610 ( .A(n1240), .B(n877), .S(n852), .Z(n726) );
  MUX21L U611 ( .A(n1239), .B(n878), .S(n852), .Z(n725) );
  MUX21L U612 ( .A(n1238), .B(n879), .S(n852), .Z(n724) );
  MUX21L U613 ( .A(n1237), .B(n880), .S(n852), .Z(n723) );
  MUX21L U614 ( .A(n1236), .B(n881), .S(n852), .Z(n722) );
  MUX21L U615 ( .A(n1235), .B(n882), .S(n852), .Z(n721) );
  MUX21L U616 ( .A(n1234), .B(n883), .S(n852), .Z(n720) );
  MUX21L U617 ( .A(n1233), .B(n884), .S(n852), .Z(n719) );
  MUX21L U618 ( .A(n1232), .B(n885), .S(n852), .Z(n718) );
  MUX21L U619 ( .A(n1231), .B(n886), .S(n852), .Z(n717) );
  MUX21L U620 ( .A(n1230), .B(n887), .S(n852), .Z(n716) );
  AN3 U621 ( .A(n2), .B(n3), .C(n845), .Z(n852) );
  MUX21L U622 ( .A(n1229), .B(n851), .S(n888), .Z(n715) );
  MUX21L U623 ( .A(n1228), .B(n853), .S(n888), .Z(n714) );
  MUX21L U624 ( .A(n1227), .B(n854), .S(n888), .Z(n713) );
  MUX21L U625 ( .A(n1226), .B(n855), .S(n888), .Z(n712) );
  MUX21L U626 ( .A(n1225), .B(n856), .S(n888), .Z(n711) );
  MUX21L U627 ( .A(n1224), .B(n857), .S(n888), .Z(n710) );
  MUX21L U628 ( .A(n1223), .B(n858), .S(n888), .Z(n709) );
  MUX21L U629 ( .A(n1222), .B(n859), .S(n888), .Z(n708) );
  MUX21L U630 ( .A(n1221), .B(n860), .S(n888), .Z(n707) );
  MUX21L U631 ( .A(n1220), .B(n861), .S(n888), .Z(n706) );
  MUX21L U632 ( .A(n1219), .B(n862), .S(n888), .Z(n705) );
  MUX21L U633 ( .A(n1218), .B(n863), .S(n888), .Z(n704) );
  MUX21L U634 ( .A(n1217), .B(n864), .S(n888), .Z(n703) );
  MUX21L U635 ( .A(n1216), .B(n865), .S(n888), .Z(n702) );
  MUX21L U636 ( .A(n1215), .B(n866), .S(n888), .Z(n701) );
  MUX21L U637 ( .A(n1214), .B(n867), .S(n888), .Z(n700) );
  MUX21L U638 ( .A(n1213), .B(n868), .S(n888), .Z(n699) );
  MUX21L U639 ( .A(n1212), .B(n869), .S(n888), .Z(n698) );
  MUX21L U640 ( .A(n1211), .B(n870), .S(n888), .Z(n697) );
  MUX21L U641 ( .A(n1210), .B(n871), .S(n888), .Z(n696) );
  MUX21L U642 ( .A(n1209), .B(n872), .S(n888), .Z(n695) );
  MUX21L U643 ( .A(n1208), .B(n873), .S(n888), .Z(n694) );
  MUX21L U644 ( .A(n1207), .B(n874), .S(n888), .Z(n693) );
  MUX21L U645 ( .A(n1206), .B(n875), .S(n888), .Z(n692) );
  MUX21L U646 ( .A(n1205), .B(n876), .S(n888), .Z(n691) );
  MUX21L U647 ( .A(n1204), .B(n877), .S(n888), .Z(n690) );
  MUX21L U648 ( .A(n1203), .B(n878), .S(n888), .Z(n689) );
  MUX21L U649 ( .A(n1202), .B(n879), .S(n888), .Z(n688) );
  MUX21L U650 ( .A(n1201), .B(n880), .S(n888), .Z(n687) );
  MUX21L U651 ( .A(n1200), .B(n881), .S(n888), .Z(n686) );
  MUX21L U652 ( .A(n1199), .B(n882), .S(n888), .Z(n685) );
  MUX21L U653 ( .A(n1198), .B(n883), .S(n888), .Z(n684) );
  MUX21L U654 ( .A(n1197), .B(n884), .S(n888), .Z(n683) );
  MUX21L U655 ( .A(n1196), .B(n885), .S(n888), .Z(n682) );
  MUX21L U656 ( .A(n1195), .B(n886), .S(n888), .Z(n681) );
  MUX21L U657 ( .A(n1194), .B(n887), .S(n888), .Z(n680) );
  AN3 U658 ( .A(wr_en), .B(n2), .C(n889), .Z(n888) );
  MUX21L U659 ( .A(n1193), .B(n851), .S(n890), .Z(n679) );
  MUX21L U660 ( .A(n1192), .B(n853), .S(n890), .Z(n678) );
  MUX21L U661 ( .A(n1191), .B(n854), .S(n890), .Z(n677) );
  MUX21L U662 ( .A(n1190), .B(n855), .S(n890), .Z(n676) );
  MUX21L U663 ( .A(n1189), .B(n856), .S(n890), .Z(n675) );
  MUX21L U664 ( .A(n1188), .B(n857), .S(n890), .Z(n674) );
  MUX21L U665 ( .A(n1187), .B(n858), .S(n890), .Z(n673) );
  MUX21L U666 ( .A(n1186), .B(n859), .S(n890), .Z(n672) );
  MUX21L U667 ( .A(n1185), .B(n860), .S(n890), .Z(n671) );
  MUX21L U668 ( .A(n1184), .B(n861), .S(n890), .Z(n670) );
  MUX21L U669 ( .A(n1183), .B(n862), .S(n890), .Z(n669) );
  MUX21L U670 ( .A(n1182), .B(n863), .S(n890), .Z(n668) );
  MUX21L U671 ( .A(n1181), .B(n864), .S(n890), .Z(n667) );
  MUX21L U672 ( .A(n1180), .B(n865), .S(n890), .Z(n666) );
  MUX21L U673 ( .A(n1179), .B(n866), .S(n890), .Z(n665) );
  MUX21L U674 ( .A(n1178), .B(n867), .S(n890), .Z(n664) );
  MUX21L U675 ( .A(n1177), .B(n868), .S(n890), .Z(n663) );
  MUX21L U676 ( .A(n1176), .B(n869), .S(n890), .Z(n662) );
  MUX21L U677 ( .A(n1175), .B(n870), .S(n890), .Z(n661) );
  MUX21L U678 ( .A(n1174), .B(n871), .S(n890), .Z(n660) );
  MUX21L U679 ( .A(n1173), .B(n872), .S(n890), .Z(n659) );
  MUX21L U680 ( .A(n1172), .B(n873), .S(n890), .Z(n658) );
  MUX21L U681 ( .A(n1171), .B(n874), .S(n890), .Z(n657) );
  MUX21L U682 ( .A(n1170), .B(n875), .S(n890), .Z(n656) );
  MUX21L U683 ( .A(n1169), .B(n876), .S(n890), .Z(n655) );
  MUX21L U684 ( .A(n1168), .B(n877), .S(n890), .Z(n654) );
  MUX21L U685 ( .A(n1167), .B(n878), .S(n890), .Z(n653) );
  MUX21L U686 ( .A(n1166), .B(n879), .S(n890), .Z(n652) );
  MUX21L U687 ( .A(n1165), .B(n880), .S(n890), .Z(n651) );
  MUX21L U688 ( .A(n1164), .B(n881), .S(n890), .Z(n650) );
  MUX21L U689 ( .A(n1163), .B(n882), .S(n890), .Z(n649) );
  MUX21L U690 ( .A(n1162), .B(n883), .S(n890), .Z(n648) );
  MUX21L U691 ( .A(n1161), .B(n884), .S(n890), .Z(n647) );
  MUX21L U692 ( .A(n1160), .B(n885), .S(n890), .Z(n646) );
  MUX21L U693 ( .A(n1159), .B(n886), .S(n890), .Z(n645) );
  MUX21L U694 ( .A(n1158), .B(n887), .S(n890), .Z(n644) );
  AN3 U695 ( .A(n2), .B(wr_ptr_1_), .C(n845), .Z(n890) );
  MUX21L U696 ( .A(n1157), .B(n851), .S(n891), .Z(n643) );
  MUX21L U697 ( .A(n1156), .B(n853), .S(n891), .Z(n642) );
  MUX21L U698 ( .A(n1155), .B(n854), .S(n891), .Z(n641) );
  MUX21L U699 ( .A(n1154), .B(n855), .S(n891), .Z(n640) );
  MUX21L U700 ( .A(n1153), .B(n856), .S(n891), .Z(n639) );
  MUX21L U701 ( .A(n1152), .B(n857), .S(n891), .Z(n638) );
  MUX21L U702 ( .A(n1151), .B(n858), .S(n891), .Z(n637) );
  MUX21L U703 ( .A(n1150), .B(n859), .S(n891), .Z(n636) );
  MUX21L U704 ( .A(n1149), .B(n860), .S(n891), .Z(n635) );
  MUX21L U705 ( .A(n1148), .B(n861), .S(n891), .Z(n634) );
  MUX21L U706 ( .A(n1147), .B(n862), .S(n891), .Z(n633) );
  MUX21L U707 ( .A(n1146), .B(n863), .S(n891), .Z(n632) );
  MUX21L U708 ( .A(n1145), .B(n864), .S(n891), .Z(n631) );
  MUX21L U709 ( .A(n1144), .B(n865), .S(n891), .Z(n630) );
  MUX21L U710 ( .A(n1143), .B(n866), .S(n891), .Z(n629) );
  MUX21L U711 ( .A(n1142), .B(n867), .S(n891), .Z(n628) );
  MUX21L U712 ( .A(n1141), .B(n868), .S(n891), .Z(n627) );
  MUX21L U713 ( .A(n1140), .B(n869), .S(n891), .Z(n626) );
  MUX21L U714 ( .A(n1139), .B(n870), .S(n891), .Z(n625) );
  MUX21L U715 ( .A(n1138), .B(n871), .S(n891), .Z(n624) );
  MUX21L U716 ( .A(n1137), .B(n872), .S(n891), .Z(n623) );
  MUX21L U717 ( .A(n1136), .B(n873), .S(n891), .Z(n622) );
  MUX21L U718 ( .A(n1135), .B(n874), .S(n891), .Z(n621) );
  MUX21L U719 ( .A(n1134), .B(n875), .S(n891), .Z(n620) );
  MUX21L U720 ( .A(n1133), .B(n876), .S(n891), .Z(n619) );
  MUX21L U721 ( .A(n1132), .B(n877), .S(n891), .Z(n618) );
  MUX21L U722 ( .A(n1131), .B(n878), .S(n891), .Z(n617) );
  MUX21L U723 ( .A(n1130), .B(n879), .S(n891), .Z(n616) );
  MUX21L U724 ( .A(n1129), .B(n880), .S(n891), .Z(n615) );
  MUX21L U725 ( .A(n1128), .B(n881), .S(n891), .Z(n614) );
  MUX21L U726 ( .A(n1127), .B(n882), .S(n891), .Z(n613) );
  MUX21L U727 ( .A(n1126), .B(n883), .S(n891), .Z(n612) );
  MUX21L U728 ( .A(n1125), .B(n884), .S(n891), .Z(n611) );
  MUX21L U729 ( .A(n1124), .B(n885), .S(n891), .Z(n610) );
  MUX21L U730 ( .A(n1123), .B(n886), .S(n891), .Z(n609) );
  MUX21L U731 ( .A(n1122), .B(n887), .S(n891), .Z(n608) );
  AN3 U732 ( .A(n2), .B(wr_en), .C(n892), .Z(n891) );
  MUX21L U733 ( .A(n1121), .B(n851), .S(n893), .Z(n607) );
  MUX21L U734 ( .A(n1120), .B(n853), .S(n893), .Z(n606) );
  MUX21L U735 ( .A(n1119), .B(n854), .S(n893), .Z(n605) );
  MUX21L U736 ( .A(n1118), .B(n855), .S(n893), .Z(n604) );
  MUX21L U737 ( .A(n1117), .B(n856), .S(n893), .Z(n603) );
  MUX21L U738 ( .A(n1116), .B(n857), .S(n893), .Z(n602) );
  MUX21L U739 ( .A(n1115), .B(n858), .S(n893), .Z(n601) );
  MUX21L U740 ( .A(n1114), .B(n859), .S(n893), .Z(n600) );
  MUX21L U741 ( .A(n1113), .B(n860), .S(n893), .Z(n599) );
  MUX21L U742 ( .A(n1112), .B(n861), .S(n893), .Z(n598) );
  MUX21L U743 ( .A(n1111), .B(n862), .S(n893), .Z(n597) );
  MUX21L U744 ( .A(n1110), .B(n863), .S(n893), .Z(n596) );
  MUX21L U745 ( .A(n1109), .B(n864), .S(n893), .Z(n595) );
  MUX21L U746 ( .A(n1108), .B(n865), .S(n893), .Z(n594) );
  MUX21L U747 ( .A(n1107), .B(n866), .S(n893), .Z(n593) );
  MUX21L U748 ( .A(n1106), .B(n867), .S(n893), .Z(n592) );
  MUX21L U749 ( .A(n1105), .B(n868), .S(n893), .Z(n591) );
  MUX21L U750 ( .A(n1104), .B(n869), .S(n893), .Z(n590) );
  MUX21L U751 ( .A(n1103), .B(n870), .S(n893), .Z(n589) );
  MUX21L U752 ( .A(n1102), .B(n871), .S(n893), .Z(n588) );
  MUX21L U753 ( .A(n1101), .B(n872), .S(n893), .Z(n587) );
  MUX21L U754 ( .A(n1100), .B(n873), .S(n893), .Z(n586) );
  MUX21L U755 ( .A(n1099), .B(n874), .S(n893), .Z(n585) );
  MUX21L U756 ( .A(n1098), .B(n875), .S(n893), .Z(n584) );
  MUX21L U757 ( .A(n1097), .B(n876), .S(n893), .Z(n583) );
  MUX21L U758 ( .A(n1096), .B(n877), .S(n893), .Z(n582) );
  MUX21L U759 ( .A(n1095), .B(n878), .S(n893), .Z(n581) );
  MUX21L U760 ( .A(n1094), .B(n879), .S(n893), .Z(n580) );
  MUX21L U761 ( .A(n1093), .B(n880), .S(n893), .Z(n579) );
  MUX21L U762 ( .A(n1092), .B(n881), .S(n893), .Z(n578) );
  MUX21L U763 ( .A(n1091), .B(n882), .S(n893), .Z(n577) );
  MUX21L U764 ( .A(n1090), .B(n883), .S(n893), .Z(n576) );
  MUX21L U765 ( .A(n1089), .B(n884), .S(n893), .Z(n575) );
  MUX21L U766 ( .A(n1088), .B(n885), .S(n893), .Z(n574) );
  MUX21L U767 ( .A(n1087), .B(n886), .S(n893), .Z(n573) );
  MUX21L U768 ( .A(n1086), .B(n887), .S(n893), .Z(n572) );
  AN3 U769 ( .A(n3), .B(wr_ptr_2_), .C(n845), .Z(n893) );
  MUX21L U770 ( .A(n1085), .B(n851), .S(n894), .Z(n571) );
  MUX21L U771 ( .A(n1084), .B(n853), .S(n894), .Z(n570) );
  MUX21L U772 ( .A(n1083), .B(n854), .S(n894), .Z(n569) );
  MUX21L U773 ( .A(n1082), .B(n855), .S(n894), .Z(n568) );
  MUX21L U774 ( .A(n1081), .B(n856), .S(n894), .Z(n567) );
  MUX21L U775 ( .A(n1080), .B(n857), .S(n894), .Z(n566) );
  MUX21L U776 ( .A(n1079), .B(n858), .S(n894), .Z(n565) );
  MUX21L U777 ( .A(n1078), .B(n859), .S(n894), .Z(n564) );
  MUX21L U778 ( .A(n1077), .B(n860), .S(n894), .Z(n563) );
  MUX21L U779 ( .A(n1076), .B(n861), .S(n894), .Z(n562) );
  MUX21L U780 ( .A(n1075), .B(n862), .S(n894), .Z(n561) );
  MUX21L U781 ( .A(n1074), .B(n863), .S(n894), .Z(n560) );
  MUX21L U782 ( .A(n1073), .B(n864), .S(n894), .Z(n559) );
  MUX21L U783 ( .A(n1072), .B(n865), .S(n894), .Z(n558) );
  MUX21L U784 ( .A(n1071), .B(n866), .S(n894), .Z(n557) );
  MUX21L U785 ( .A(n1070), .B(n867), .S(n894), .Z(n556) );
  MUX21L U786 ( .A(n1069), .B(n868), .S(n894), .Z(n555) );
  MUX21L U787 ( .A(n1068), .B(n869), .S(n894), .Z(n554) );
  MUX21L U788 ( .A(n1067), .B(n870), .S(n894), .Z(n553) );
  MUX21L U789 ( .A(n1066), .B(n871), .S(n894), .Z(n552) );
  MUX21L U790 ( .A(n1065), .B(n872), .S(n894), .Z(n551) );
  MUX21L U791 ( .A(n1064), .B(n873), .S(n894), .Z(n550) );
  MUX21L U792 ( .A(n1063), .B(n874), .S(n894), .Z(n549) );
  MUX21L U793 ( .A(n1062), .B(n875), .S(n894), .Z(n548) );
  MUX21L U794 ( .A(n1061), .B(n876), .S(n894), .Z(n547) );
  MUX21L U795 ( .A(n1060), .B(n877), .S(n894), .Z(n546) );
  MUX21L U796 ( .A(n1059), .B(n878), .S(n894), .Z(n545) );
  MUX21L U797 ( .A(n1058), .B(n879), .S(n894), .Z(n544) );
  MUX21L U798 ( .A(n1057), .B(n880), .S(n894), .Z(n543) );
  MUX21L U799 ( .A(n1056), .B(n881), .S(n894), .Z(n542) );
  MUX21L U800 ( .A(n1055), .B(n882), .S(n894), .Z(n541) );
  MUX21L U801 ( .A(n1054), .B(n883), .S(n894), .Z(n540) );
  MUX21L U802 ( .A(n1053), .B(n884), .S(n894), .Z(n539) );
  MUX21L U803 ( .A(n1052), .B(n885), .S(n894), .Z(n538) );
  MUX21L U804 ( .A(n1051), .B(n886), .S(n894), .Z(n537) );
  MUX21L U805 ( .A(n1050), .B(n887), .S(n894), .Z(n536) );
  AN3 U806 ( .A(wr_ptr_2_), .B(wr_en), .C(n889), .Z(n894) );
  MUX21L U807 ( .A(n1049), .B(n851), .S(n895), .Z(n535) );
  MUX21L U808 ( .A(n1048), .B(n853), .S(n895), .Z(n534) );
  MUX21L U809 ( .A(n1047), .B(n854), .S(n895), .Z(n533) );
  MUX21L U810 ( .A(n1046), .B(n855), .S(n895), .Z(n532) );
  MUX21L U811 ( .A(n1045), .B(n856), .S(n895), .Z(n531) );
  MUX21L U812 ( .A(n1044), .B(n857), .S(n895), .Z(n530) );
  MUX21L U813 ( .A(n1043), .B(n858), .S(n895), .Z(n529) );
  MUX21L U814 ( .A(n1042), .B(n859), .S(n895), .Z(n528) );
  MUX21L U815 ( .A(n1041), .B(n860), .S(n895), .Z(n527) );
  MUX21L U816 ( .A(n1040), .B(n861), .S(n895), .Z(n526) );
  MUX21L U817 ( .A(n1039), .B(n862), .S(n895), .Z(n525) );
  MUX21L U818 ( .A(n1038), .B(n863), .S(n895), .Z(n524) );
  MUX21L U819 ( .A(n1037), .B(n864), .S(n895), .Z(n523) );
  MUX21L U820 ( .A(n1036), .B(n865), .S(n895), .Z(n522) );
  MUX21L U821 ( .A(n1035), .B(n866), .S(n895), .Z(n521) );
  MUX21L U822 ( .A(n1034), .B(n867), .S(n895), .Z(n520) );
  MUX21L U823 ( .A(n1033), .B(n868), .S(n895), .Z(n519) );
  MUX21L U824 ( .A(n1032), .B(n869), .S(n895), .Z(n518) );
  MUX21L U825 ( .A(n1031), .B(n870), .S(n895), .Z(n517) );
  MUX21L U826 ( .A(n1030), .B(n871), .S(n895), .Z(n516) );
  MUX21L U827 ( .A(n1029), .B(n872), .S(n895), .Z(n515) );
  MUX21L U828 ( .A(n1028), .B(n873), .S(n895), .Z(n514) );
  MUX21L U829 ( .A(n1027), .B(n874), .S(n895), .Z(n513) );
  MUX21L U830 ( .A(n1026), .B(n875), .S(n895), .Z(n512) );
  MUX21L U831 ( .A(n1025), .B(n876), .S(n895), .Z(n511) );
  MUX21L U832 ( .A(n1024), .B(n877), .S(n895), .Z(n510) );
  MUX21L U833 ( .A(n1023), .B(n878), .S(n895), .Z(n509) );
  MUX21L U834 ( .A(n1022), .B(n879), .S(n895), .Z(n508) );
  MUX21L U835 ( .A(n1021), .B(n880), .S(n895), .Z(n507) );
  MUX21L U836 ( .A(n1020), .B(n881), .S(n895), .Z(n506) );
  MUX21L U837 ( .A(n1019), .B(n882), .S(n895), .Z(n505) );
  MUX21L U838 ( .A(n1018), .B(n883), .S(n895), .Z(n504) );
  MUX21L U839 ( .A(n1017), .B(n884), .S(n895), .Z(n503) );
  MUX21L U840 ( .A(n1016), .B(n885), .S(n895), .Z(n502) );
  MUX21L U841 ( .A(n1015), .B(n886), .S(n895), .Z(n501) );
  MUX21L U842 ( .A(n1014), .B(n887), .S(n895), .Z(n500) );
  AN3 U843 ( .A(wr_ptr_1_), .B(wr_ptr_2_), .C(n845), .Z(n895) );
  MUX21L U844 ( .A(n1013), .B(n851), .S(n896), .Z(n499) );
  IV U845 ( .A(wr_data[0]), .Z(n851) );
  MUX21L U846 ( .A(n1012), .B(n853), .S(n896), .Z(n498) );
  IV U847 ( .A(wr_data[35]), .Z(n853) );
  MUX21L U848 ( .A(n1011), .B(n854), .S(n896), .Z(n497) );
  IV U849 ( .A(wr_data[34]), .Z(n854) );
  MUX21L U850 ( .A(n1010), .B(n855), .S(n896), .Z(n496) );
  IV U851 ( .A(wr_data[33]), .Z(n855) );
  MUX21L U852 ( .A(n1009), .B(n856), .S(n896), .Z(n495) );
  IV U853 ( .A(wr_data[32]), .Z(n856) );
  MUX21L U854 ( .A(n1008), .B(n857), .S(n896), .Z(n494) );
  IV U855 ( .A(wr_data[31]), .Z(n857) );
  MUX21L U856 ( .A(n1007), .B(n858), .S(n896), .Z(n493) );
  IV U857 ( .A(wr_data[30]), .Z(n858) );
  MUX21L U858 ( .A(n1006), .B(n859), .S(n896), .Z(n492) );
  IV U859 ( .A(wr_data[29]), .Z(n859) );
  MUX21L U860 ( .A(n1005), .B(n860), .S(n896), .Z(n491) );
  IV U861 ( .A(wr_data[28]), .Z(n860) );
  MUX21L U862 ( .A(n1004), .B(n861), .S(n896), .Z(n490) );
  IV U863 ( .A(wr_data[27]), .Z(n861) );
  MUX21L U864 ( .A(n1003), .B(n862), .S(n896), .Z(n489) );
  IV U865 ( .A(wr_data[26]), .Z(n862) );
  MUX21L U866 ( .A(n1002), .B(n863), .S(n896), .Z(n488) );
  IV U867 ( .A(wr_data[25]), .Z(n863) );
  MUX21L U868 ( .A(n1001), .B(n864), .S(n896), .Z(n487) );
  IV U869 ( .A(wr_data[24]), .Z(n864) );
  MUX21L U870 ( .A(n1000), .B(n865), .S(n896), .Z(n486) );
  IV U871 ( .A(wr_data[23]), .Z(n865) );
  MUX21L U872 ( .A(n999), .B(n866), .S(n896), .Z(n485) );
  IV U873 ( .A(wr_data[22]), .Z(n866) );
  MUX21L U874 ( .A(n998), .B(n867), .S(n896), .Z(n484) );
  IV U875 ( .A(wr_data[21]), .Z(n867) );
  MUX21L U876 ( .A(n997), .B(n868), .S(n896), .Z(n483) );
  IV U877 ( .A(wr_data[20]), .Z(n868) );
  MUX21L U878 ( .A(n996), .B(n869), .S(n896), .Z(n482) );
  IV U879 ( .A(wr_data[19]), .Z(n869) );
  MUX21L U880 ( .A(n995), .B(n870), .S(n896), .Z(n481) );
  IV U881 ( .A(wr_data[18]), .Z(n870) );
  MUX21L U882 ( .A(n994), .B(n871), .S(n896), .Z(n480) );
  IV U883 ( .A(wr_data[17]), .Z(n871) );
  MUX21L U884 ( .A(n993), .B(n872), .S(n896), .Z(n479) );
  IV U885 ( .A(wr_data[16]), .Z(n872) );
  MUX21L U886 ( .A(n992), .B(n873), .S(n896), .Z(n478) );
  IV U887 ( .A(wr_data[15]), .Z(n873) );
  MUX21L U888 ( .A(n991), .B(n874), .S(n896), .Z(n477) );
  IV U889 ( .A(wr_data[14]), .Z(n874) );
  MUX21L U890 ( .A(n990), .B(n875), .S(n896), .Z(n476) );
  IV U891 ( .A(wr_data[13]), .Z(n875) );
  MUX21L U892 ( .A(n989), .B(n876), .S(n896), .Z(n475) );
  IV U893 ( .A(wr_data[12]), .Z(n876) );
  MUX21L U894 ( .A(n988), .B(n877), .S(n896), .Z(n474) );
  IV U895 ( .A(wr_data[11]), .Z(n877) );
  MUX21L U896 ( .A(n987), .B(n878), .S(n896), .Z(n473) );
  IV U897 ( .A(wr_data[10]), .Z(n878) );
  MUX21L U898 ( .A(n986), .B(n879), .S(n896), .Z(n472) );
  IV U899 ( .A(wr_data[9]), .Z(n879) );
  MUX21L U900 ( .A(n985), .B(n880), .S(n896), .Z(n471) );
  IV U901 ( .A(wr_data[8]), .Z(n880) );
  MUX21L U902 ( .A(n984), .B(n881), .S(n896), .Z(n470) );
  IV U903 ( .A(wr_data[7]), .Z(n881) );
  MUX21L U904 ( .A(n983), .B(n882), .S(n896), .Z(n469) );
  IV U905 ( .A(wr_data[6]), .Z(n882) );
  MUX21L U906 ( .A(n982), .B(n883), .S(n896), .Z(n468) );
  IV U907 ( .A(wr_data[5]), .Z(n883) );
  MUX21L U908 ( .A(n981), .B(n884), .S(n896), .Z(n467) );
  IV U909 ( .A(wr_data[4]), .Z(n884) );
  MUX21L U910 ( .A(n980), .B(n885), .S(n896), .Z(n466) );
  IV U911 ( .A(wr_data[3]), .Z(n885) );
  MUX21L U912 ( .A(n979), .B(n886), .S(n896), .Z(n465) );
  IV U913 ( .A(wr_data[2]), .Z(n886) );
  MUX21L U914 ( .A(n978), .B(n887), .S(n896), .Z(n464) );
  NR2 U915 ( .A(n897), .B(n847), .Z(n896) );
  IV U916 ( .A(wr_data[1]), .Z(n887) );
  IV U917 ( .A(n898), .Z(n463) );
  AO6 U918 ( .A(n847), .B(test_so7), .C(n899), .Z(n898) );
  AO7 U919 ( .A(wr_en), .B(n977), .C(n900), .Z(n462) );
  AO2 U920 ( .A(n899), .B(n901), .C(n850), .D(n902), .Z(n900) );
  AO7 U921 ( .A(wr_en), .B(n976), .C(n903), .Z(n461) );
  IV U922 ( .A(n899), .Z(n903) );
  NR2 U923 ( .A(n847), .B(n902), .Z(n899) );
  EO U924 ( .A(test_so7), .B(n897), .Z(n902) );
  AO7 U925 ( .A(wr_en), .B(n975), .C(n904), .Z(n460) );
  AO2 U926 ( .A(n848), .B(n1242), .C(n905), .D(n845), .Z(n904) );
  NR2 U927 ( .A(n847), .B(n1242), .Z(n845) );
  AO7 U928 ( .A(wr_en), .B(n974), .C(n906), .Z(n459) );
  AO2 U929 ( .A(n905), .B(n850), .C(n848), .D(n901), .Z(n906) );
  NR2 U930 ( .A(n847), .B(n905), .Z(n848) );
  NR2 U931 ( .A(n901), .B(n847), .Z(n850) );
  AO7 U932 ( .A(wr_ptr_2_), .B(n892), .C(n897), .Z(n901) );
  ND2 U933 ( .A(n892), .B(wr_ptr_2_), .Z(n897) );
  NR2 U934 ( .A(n3), .B(n1), .Z(n892) );
  AO6 U935 ( .A(n1), .B(wr_ptr_1_), .C(n889), .Z(n905) );
  NR2 U936 ( .A(n1), .B(wr_ptr_1_), .Z(n889) );
  AO4 U937 ( .A(n907), .B(n847), .C(n972), .D(n908), .Z(n458) );
  IV U938 ( .A(wr_en), .Z(n847) );
  NR2 U939 ( .A(afull), .B(full), .Z(n907) );
  NR2 U940 ( .A(n909), .B(n910), .Z(empty) );
  EN U941 ( .A(n911), .B(N69), .Z(n909) );
  AN4 U942 ( .A(n908), .B(n912), .C(n913), .D(n914), .Z(afull) );
  AO7 U943 ( .A(n1), .B(n915), .C(n916), .Z(n914) );
  EN U944 ( .A(n917), .B(n918), .Z(n913) );
  EN U945 ( .A(wr_ptr_1_), .B(n916), .Z(n918) );
  EO U946 ( .A(n919), .B(n920), .Z(n912) );
  EN U947 ( .A(wr_ptr_2_), .B(n921), .Z(n920) );
  AO5 U948 ( .A(n922), .B(n923), .C(n3), .Z(n921) );
  EO U949 ( .A(sync_rd_ptr_1[1]), .B(n919), .Z(n923) );
  AN2 U950 ( .A(n1), .B(n915), .Z(n922) );
  EO U951 ( .A(n924), .B(n925), .Z(n908) );
  EO U952 ( .A(test_so7), .B(sync_rd_ptr_1[3]), .Z(n925) );
  AO5 U953 ( .A(n926), .B(n927), .C(n2), .Z(n924) );
  EO U954 ( .A(sync_rd_ptr_1[3]), .B(sync_rd_ptr_1[2]), .Z(n927) );
  AO2 U955 ( .A(wr_ptr_1_), .B(n928), .C(n917), .D(n916), .Z(n926) );
  OR2 U956 ( .A(n916), .B(n917), .Z(n928) );
  ND2 U957 ( .A(n915), .B(n1), .Z(n916) );
  EN U958 ( .A(n917), .B(sync_rd_ptr_1[0]), .Z(n915) );
  EN U959 ( .A(n919), .B(sync_rd_ptr_1[1]), .Z(n917) );
  EN U960 ( .A(n973), .B(sync_rd_ptr_1[3]), .Z(n919) );
  NR2 U961 ( .A(n910), .B(n929), .Z(aempty) );
  EN U962 ( .A(n970), .B(n911), .Z(n929) );
  AO3 U963 ( .A(n930), .B(n931), .C(n932), .D(n933), .Z(n910) );
  MUX21L U964 ( .A(n934), .B(n935), .S(n936), .Z(n933) );
  AN3 U965 ( .A(n937), .B(N69), .C(n911), .Z(n936) );
  AN2 U966 ( .A(n938), .B(n931), .Z(n935) );
  AO7 U967 ( .A(n360), .B(n939), .C(n938), .Z(n934) );
  ND2 U968 ( .A(n360), .B(n939), .Z(n938) );
  EO U969 ( .A(n937), .B(n940), .Z(n932) );
  AO2 U970 ( .A(n969), .B(n941), .C(n911), .D(n837), .Z(n940) );
  NR2 U971 ( .A(n969), .B(n970), .Z(n837) );
  ND2 U972 ( .A(n911), .B(N69), .Z(n941) );
  EO U973 ( .A(n937), .B(sync_wr_ptr_1_0_), .Z(n911) );
  EN U974 ( .A(n939), .B(sync_wr_ptr_1_1_), .Z(n937) );
  EO U975 ( .A(n4), .B(test_so8), .Z(n931) );
  NR2 U976 ( .A(n360), .B(n939), .Z(n930) );
  EN U977 ( .A(n971), .B(test_so8), .Z(n939) );
endmodule
