module sdrc_req_gen_SDR_DW16_SDR_BW2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [24:1] carry;

  FA1A U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA1A U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA1A U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA1A U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA1A U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA1A U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  EO U1 ( .A(A[11]), .B(carry[11]), .Z(SUM[11]) );
  EO U2 ( .A(A[10]), .B(carry[10]), .Z(SUM[10]) );
  EO U3 ( .A(A[9]), .B(carry[9]), .Z(SUM[9]) );
  EO U4 ( .A(A[8]), .B(carry[8]), .Z(SUM[8]) );
  EO U5 ( .A(A[7]), .B(carry[7]), .Z(SUM[7]) );
  EO U6 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
  EN U7 ( .A(A[25]), .B(n1), .Z(SUM[25]) );
  ND2 U8 ( .A(A[24]), .B(carry[24]), .Z(n1) );
  EO U9 ( .A(A[24]), .B(carry[24]), .Z(SUM[24]) );
  EO U10 ( .A(A[23]), .B(carry[23]), .Z(SUM[23]) );
  EO U11 ( .A(A[22]), .B(carry[22]), .Z(SUM[22]) );
  EO U12 ( .A(A[21]), .B(carry[21]), .Z(SUM[21]) );
  EO U13 ( .A(A[20]), .B(carry[20]), .Z(SUM[20]) );
  EO U14 ( .A(A[19]), .B(carry[19]), .Z(SUM[19]) );
  EO U15 ( .A(A[18]), .B(carry[18]), .Z(SUM[18]) );
  EO U16 ( .A(A[17]), .B(carry[17]), .Z(SUM[17]) );
  EO U17 ( .A(A[16]), .B(carry[16]), .Z(SUM[16]) );
  EO U18 ( .A(A[15]), .B(carry[15]), .Z(SUM[15]) );
  EO U19 ( .A(A[14]), .B(carry[14]), .Z(SUM[14]) );
  EO U20 ( .A(A[13]), .B(carry[13]), .Z(SUM[13]) );
  EO U21 ( .A(A[12]), .B(carry[12]), .Z(SUM[12]) );
  AN2P U22 ( .A(A[23]), .B(carry[23]), .Z(carry[24]) );
  AN2P U23 ( .A(A[22]), .B(carry[22]), .Z(carry[23]) );
  AN2P U24 ( .A(A[21]), .B(carry[21]), .Z(carry[22]) );
  AN2P U25 ( .A(A[20]), .B(carry[20]), .Z(carry[21]) );
  AN2P U26 ( .A(A[19]), .B(carry[19]), .Z(carry[20]) );
  AN2P U27 ( .A(A[18]), .B(carry[18]), .Z(carry[19]) );
  AN2P U28 ( .A(A[17]), .B(carry[17]), .Z(carry[18]) );
  AN2P U29 ( .A(A[16]), .B(carry[16]), .Z(carry[17]) );
  AN2P U30 ( .A(A[15]), .B(carry[15]), .Z(carry[16]) );
  AN2P U31 ( .A(A[14]), .B(carry[14]), .Z(carry[15]) );
  AN2P U32 ( .A(A[13]), .B(carry[13]), .Z(carry[14]) );
  AN2P U33 ( .A(A[12]), .B(carry[12]), .Z(carry[13]) );
  AN2P U34 ( .A(A[11]), .B(carry[11]), .Z(carry[12]) );
  AN2P U35 ( .A(A[10]), .B(carry[10]), .Z(carry[11]) );
  AN2P U36 ( .A(A[9]), .B(carry[9]), .Z(carry[10]) );
  AN2P U37 ( .A(A[8]), .B(carry[8]), .Z(carry[9]) );
  AN2P U38 ( .A(A[7]), .B(carry[7]), .Z(carry[8]) );
  AN2P U39 ( .A(A[0]), .B(B[0]), .Z(carry[1]) );
endmodule
