module async_fifo_36_4_0_0_test_1 ( wr_clk, wr_reset_n, wr_en, wr_data, full, 
        afull, rd_clk, rd_reset_n, rd_en, empty, aempty, rd_data, test_si6, 
        test_si5, test_si4, test_si3, test_si2, test_si1, test_so5, test_so4, 
        test_so3, test_so2, test_so1, test_se );
  input [35:0] wr_data;
  output [35:0] rd_data;
  input wr_clk, wr_reset_n, wr_en, rd_clk, rd_reset_n, rd_en, test_si6,
         test_si5, test_si4, test_si3, test_si2, test_si1, test_se;
  output full, afull, empty, aempty, test_so5, test_so4, test_so3, test_so2,
         test_so1;
  wire   N45, N46, mem_3__35_, mem_3__34_, mem_3__33_, mem_3__32_, mem_3__31_,
         mem_3__29_, mem_3__28_, mem_3__27_, mem_3__26_, mem_3__25_,
         mem_3__24_, mem_3__23_, mem_3__22_, mem_3__21_, mem_3__20_,
         mem_3__19_, mem_3__18_, mem_3__17_, mem_3__16_, mem_3__15_,
         mem_3__14_, mem_3__13_, mem_3__12_, mem_3__11_, mem_3__10_, mem_3__9_,
         mem_3__8_, mem_3__7_, mem_3__6_, mem_3__5_, mem_3__4_, mem_3__3_,
         mem_3__2_, mem_3__1_, mem_3__0_, mem_2__35_, mem_2__34_, mem_2__33_,
         mem_2__32_, mem_2__31_, mem_2__30_, mem_2__29_, mem_2__28_,
         mem_2__27_, mem_2__26_, mem_2__25_, mem_2__24_, mem_2__23_,
         mem_2__22_, mem_2__21_, mem_2__20_, mem_2__19_, mem_2__17_,
         mem_2__16_, mem_2__15_, mem_2__14_, mem_2__13_, mem_2__12_,
         mem_2__11_, mem_2__10_, mem_2__9_, mem_2__8_, mem_2__7_, mem_2__6_,
         mem_2__5_, mem_2__4_, mem_2__3_, mem_2__2_, mem_2__1_, mem_2__0_,
         mem_1__35_, mem_1__34_, mem_1__33_, mem_1__32_, mem_1__31_,
         mem_1__30_, mem_1__29_, mem_1__28_, mem_1__27_, mem_1__26_,
         mem_1__25_, mem_1__24_, mem_1__23_, mem_1__22_, mem_1__21_,
         mem_1__20_, mem_1__19_, mem_1__18_, mem_1__17_, mem_1__16_,
         mem_1__15_, mem_1__14_, mem_1__13_, mem_1__12_, mem_1__11_,
         mem_1__10_, mem_1__9_, mem_1__8_, mem_1__7_, mem_1__5_, mem_1__4_,
         mem_1__3_, mem_1__2_, mem_1__1_, mem_1__0_, mem_0__35_, mem_0__34_,
         mem_0__33_, mem_0__32_, mem_0__31_, mem_0__30_, mem_0__29_,
         mem_0__28_, mem_0__27_, mem_0__26_, mem_0__25_, mem_0__24_,
         mem_0__23_, mem_0__22_, mem_0__21_, mem_0__20_, mem_0__19_,
         mem_0__18_, mem_0__17_, mem_0__16_, mem_0__15_, mem_0__14_,
         mem_0__13_, mem_0__12_, mem_0__11_, mem_0__10_, mem_0__9_, mem_0__8_,
         mem_0__7_, mem_0__6_, mem_0__5_, mem_0__4_, mem_0__3_, mem_0__2_,
         mem_0__1_, mem_0__0_, sync_wr_ptr_1_0_, n246, n248, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n247, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n711, n712, n713, n714, n716;
  wire   [1:0] wr_ptr;
  wire   [2:0] grey_wr_ptr;
  wire   [2:0] grey_rd_ptr_dly;
  wire   [2:0] sync_rd_ptr_1;
  wire   [2:0] sync_rd_ptr_0;
  wire   [35:0] rd_data_c;
  wire   [2:0] sync_wr_ptr_0;

  FD2S sync_wr_ptr_1_reg_1_ ( .D(sync_wr_ptr_0[1]), .TI(sync_wr_ptr_1_0_), 
        .TE(test_se), .CP(n5), .CD(rd_reset_n), .Q(n716), .QN(n713) );
  FD1S mem_reg_3__35_ ( .D(n373), .TI(mem_3__34_), .TE(test_se), .CP(n17), .Q(
        mem_3__35_), .QN(n598) );
  FD1S mem_reg_3__34_ ( .D(n372), .TI(mem_3__33_), .TE(test_se), .CP(n17), .Q(
        mem_3__34_), .QN(n597) );
  FD1S mem_reg_3__33_ ( .D(n371), .TI(mem_3__32_), .TE(test_se), .CP(n17), .Q(
        mem_3__33_), .QN(n596) );
  FD1S mem_reg_3__32_ ( .D(n370), .TI(mem_3__31_), .TE(test_se), .CP(n17), .Q(
        mem_3__32_), .QN(n595) );
  FD1S mem_reg_3__31_ ( .D(n369), .TI(test_si4), .TE(test_se), .CP(n17), .Q(
        mem_3__31_), .QN(n594) );
  FD1S mem_reg_3__30_ ( .D(n368), .TI(mem_3__29_), .TE(test_se), .CP(n16), .Q(
        test_so3), .QN(n593) );
  FD1S mem_reg_3__29_ ( .D(n367), .TI(mem_3__28_), .TE(test_se), .CP(n16), .Q(
        mem_3__29_), .QN(n592) );
  FD1S mem_reg_3__28_ ( .D(n366), .TI(mem_3__27_), .TE(test_se), .CP(n16), .Q(
        mem_3__28_), .QN(n591) );
  FD1S mem_reg_3__27_ ( .D(n365), .TI(mem_3__26_), .TE(test_se), .CP(n16), .Q(
        mem_3__27_), .QN(n590) );
  FD1S mem_reg_3__26_ ( .D(n364), .TI(mem_3__25_), .TE(test_se), .CP(n16), .Q(
        mem_3__26_), .QN(n589) );
  FD1S mem_reg_3__25_ ( .D(n363), .TI(mem_3__24_), .TE(test_se), .CP(n16), .Q(
        mem_3__25_), .QN(n588) );
  FD1S mem_reg_3__24_ ( .D(n362), .TI(mem_3__23_), .TE(test_se), .CP(n16), .Q(
        mem_3__24_), .QN(n587) );
  FD1S mem_reg_3__23_ ( .D(n361), .TI(mem_3__22_), .TE(test_se), .CP(n16), .Q(
        mem_3__23_), .QN(n586) );
  FD1S mem_reg_3__22_ ( .D(n360), .TI(mem_3__21_), .TE(test_se), .CP(n16), .Q(
        mem_3__22_), .QN(n585) );
  FD1S mem_reg_3__21_ ( .D(n359), .TI(mem_3__20_), .TE(test_se), .CP(n16), .Q(
        mem_3__21_), .QN(n584) );
  FD1S mem_reg_3__20_ ( .D(n358), .TI(mem_3__19_), .TE(test_se), .CP(n16), .Q(
        mem_3__20_), .QN(n583) );
  FD1S mem_reg_3__19_ ( .D(n357), .TI(mem_3__18_), .TE(test_se), .CP(n16), .Q(
        mem_3__19_), .QN(n582) );
  FD1S mem_reg_3__18_ ( .D(n356), .TI(mem_3__17_), .TE(test_se), .CP(n15), .Q(
        mem_3__18_), .QN(n581) );
  FD1S mem_reg_3__17_ ( .D(n355), .TI(mem_3__16_), .TE(test_se), .CP(n15), .Q(
        mem_3__17_), .QN(n580) );
  FD1S mem_reg_3__16_ ( .D(n354), .TI(mem_3__15_), .TE(test_se), .CP(n15), .Q(
        mem_3__16_), .QN(n579) );
  FD1S mem_reg_3__15_ ( .D(n353), .TI(mem_3__14_), .TE(test_se), .CP(n15), .Q(
        mem_3__15_), .QN(n578) );
  FD1S mem_reg_3__14_ ( .D(n352), .TI(mem_3__13_), .TE(test_se), .CP(n15), .Q(
        mem_3__14_), .QN(n577) );
  FD1S mem_reg_3__13_ ( .D(n351), .TI(mem_3__12_), .TE(test_se), .CP(n15), .Q(
        mem_3__13_), .QN(n576) );
  FD1S mem_reg_3__12_ ( .D(n350), .TI(mem_3__11_), .TE(test_se), .CP(n15), .Q(
        mem_3__12_), .QN(n575) );
  FD1S mem_reg_3__11_ ( .D(n349), .TI(mem_3__10_), .TE(test_se), .CP(n15), .Q(
        mem_3__11_), .QN(n574) );
  FD1S mem_reg_3__10_ ( .D(n348), .TI(mem_3__9_), .TE(test_se), .CP(n15), .Q(
        mem_3__10_), .QN(n573) );
  FD1S mem_reg_3__9_ ( .D(n347), .TI(mem_3__8_), .TE(test_se), .CP(n15), .Q(
        mem_3__9_), .QN(n572) );
  FD1S mem_reg_3__8_ ( .D(n346), .TI(mem_3__7_), .TE(test_se), .CP(n15), .Q(
        mem_3__8_), .QN(n571) );
  FD1S mem_reg_3__7_ ( .D(n345), .TI(mem_3__6_), .TE(test_se), .CP(n15), .Q(
        mem_3__7_), .QN(n570) );
  FD1S mem_reg_3__6_ ( .D(n344), .TI(mem_3__5_), .TE(test_se), .CP(n14), .Q(
        mem_3__6_), .QN(n569) );
  FD1S mem_reg_3__5_ ( .D(n343), .TI(mem_3__4_), .TE(test_se), .CP(n14), .Q(
        mem_3__5_), .QN(n568) );
  FD1S mem_reg_3__4_ ( .D(n342), .TI(mem_3__3_), .TE(test_se), .CP(n14), .Q(
        mem_3__4_), .QN(n567) );
  FD1S mem_reg_3__3_ ( .D(n341), .TI(mem_3__2_), .TE(test_se), .CP(n14), .Q(
        mem_3__3_), .QN(n566) );
  FD1S mem_reg_3__2_ ( .D(n340), .TI(mem_3__1_), .TE(test_se), .CP(n14), .Q(
        mem_3__2_), .QN(n565) );
  FD1S mem_reg_3__1_ ( .D(n339), .TI(mem_3__0_), .TE(test_se), .CP(n14), .Q(
        mem_3__1_), .QN(n564) );
  FD1S mem_reg_3__0_ ( .D(n374), .TI(mem_2__35_), .TE(test_se), .CP(n17), .Q(
        mem_3__0_), .QN(n599) );
  FD1S mem_reg_2__35_ ( .D(n409), .TI(mem_2__34_), .TE(test_se), .CP(n20), .Q(
        mem_2__35_), .QN(n634) );
  FD1S mem_reg_2__34_ ( .D(n408), .TI(mem_2__33_), .TE(test_se), .CP(n20), .Q(
        mem_2__34_), .QN(n633) );
  FD1S mem_reg_2__33_ ( .D(n407), .TI(mem_2__32_), .TE(test_se), .CP(n20), .Q(
        mem_2__33_), .QN(n632) );
  FD1S mem_reg_2__32_ ( .D(n406), .TI(mem_2__31_), .TE(test_se), .CP(n20), .Q(
        mem_2__32_), .QN(n631) );
  FD1S mem_reg_2__31_ ( .D(n405), .TI(mem_2__30_), .TE(test_se), .CP(n20), .Q(
        mem_2__31_), .QN(n630) );
  FD1S mem_reg_2__30_ ( .D(n404), .TI(mem_2__29_), .TE(test_se), .CP(n19), .Q(
        mem_2__30_), .QN(n629) );
  FD1S mem_reg_2__29_ ( .D(n403), .TI(mem_2__28_), .TE(test_se), .CP(n19), .Q(
        mem_2__29_), .QN(n628) );
  FD1S mem_reg_2__28_ ( .D(n402), .TI(mem_2__27_), .TE(test_se), .CP(n19), .Q(
        mem_2__28_), .QN(n627) );
  FD1S mem_reg_2__27_ ( .D(n401), .TI(mem_2__26_), .TE(test_se), .CP(n19), .Q(
        mem_2__27_), .QN(n626) );
  FD1S mem_reg_2__26_ ( .D(n400), .TI(mem_2__25_), .TE(test_se), .CP(n19), .Q(
        mem_2__26_), .QN(n625) );
  FD1S mem_reg_2__25_ ( .D(n399), .TI(mem_2__24_), .TE(test_se), .CP(n19), .Q(
        mem_2__25_), .QN(n624) );
  FD1S mem_reg_2__24_ ( .D(n398), .TI(mem_2__23_), .TE(test_se), .CP(n19), .Q(
        mem_2__24_), .QN(n623) );
  FD1S mem_reg_2__23_ ( .D(n397), .TI(mem_2__22_), .TE(test_se), .CP(n19), .Q(
        mem_2__23_), .QN(n622) );
  FD1S mem_reg_2__22_ ( .D(n396), .TI(mem_2__21_), .TE(test_se), .CP(n19), .Q(
        mem_2__22_), .QN(n621) );
  FD1S mem_reg_2__21_ ( .D(n395), .TI(mem_2__20_), .TE(test_se), .CP(n19), .Q(
        mem_2__21_), .QN(n620) );
  FD1S mem_reg_2__20_ ( .D(n394), .TI(mem_2__19_), .TE(test_se), .CP(n19), .Q(
        mem_2__20_), .QN(n619) );
  FD1S mem_reg_2__19_ ( .D(n393), .TI(test_si3), .TE(test_se), .CP(n19), .Q(
        mem_2__19_), .QN(n618) );
  FD1S mem_reg_2__18_ ( .D(n392), .TI(mem_2__17_), .TE(test_se), .CP(n18), .Q(
        test_so2), .QN(n617) );
  FD1S mem_reg_2__17_ ( .D(n391), .TI(mem_2__16_), .TE(test_se), .CP(n18), .Q(
        mem_2__17_), .QN(n616) );
  FD1S mem_reg_2__16_ ( .D(n390), .TI(mem_2__15_), .TE(test_se), .CP(n18), .Q(
        mem_2__16_), .QN(n615) );
  FD1S mem_reg_2__15_ ( .D(n389), .TI(mem_2__14_), .TE(test_se), .CP(n18), .Q(
        mem_2__15_), .QN(n614) );
  FD1S mem_reg_2__14_ ( .D(n388), .TI(mem_2__13_), .TE(test_se), .CP(n18), .Q(
        mem_2__14_), .QN(n613) );
  FD1S mem_reg_2__13_ ( .D(n387), .TI(mem_2__12_), .TE(test_se), .CP(n18), .Q(
        mem_2__13_), .QN(n612) );
  FD1S mem_reg_2__12_ ( .D(n386), .TI(mem_2__11_), .TE(test_se), .CP(n18), .Q(
        mem_2__12_), .QN(n611) );
  FD1S mem_reg_2__11_ ( .D(n385), .TI(mem_2__10_), .TE(test_se), .CP(n18), .Q(
        mem_2__11_), .QN(n610) );
  FD1S mem_reg_2__10_ ( .D(n384), .TI(mem_2__9_), .TE(test_se), .CP(n18), .Q(
        mem_2__10_), .QN(n609) );
  FD1S mem_reg_2__9_ ( .D(n383), .TI(mem_2__8_), .TE(test_se), .CP(n18), .Q(
        mem_2__9_), .QN(n608) );
  FD1S mem_reg_2__8_ ( .D(n382), .TI(mem_2__7_), .TE(test_se), .CP(n18), .Q(
        mem_2__8_), .QN(n607) );
  FD1S mem_reg_2__7_ ( .D(n381), .TI(mem_2__6_), .TE(test_se), .CP(n18), .Q(
        mem_2__7_), .QN(n606) );
  FD1S mem_reg_2__6_ ( .D(n380), .TI(mem_2__5_), .TE(test_se), .CP(n17), .Q(
        mem_2__6_), .QN(n605) );
  FD1S mem_reg_2__5_ ( .D(n379), .TI(mem_2__4_), .TE(test_se), .CP(n17), .Q(
        mem_2__5_), .QN(n604) );
  FD1S mem_reg_2__4_ ( .D(n378), .TI(mem_2__3_), .TE(test_se), .CP(n17), .Q(
        mem_2__4_), .QN(n603) );
  FD1S mem_reg_2__3_ ( .D(n377), .TI(mem_2__2_), .TE(test_se), .CP(n17), .Q(
        mem_2__3_), .QN(n602) );
  FD1S mem_reg_2__2_ ( .D(n376), .TI(mem_2__1_), .TE(test_se), .CP(n17), .Q(
        mem_2__2_), .QN(n601) );
  FD1S mem_reg_2__1_ ( .D(n375), .TI(mem_2__0_), .TE(test_se), .CP(n17), .Q(
        mem_2__1_), .QN(n600) );
  FD1S mem_reg_2__0_ ( .D(n410), .TI(mem_1__35_), .TE(test_se), .CP(n20), .Q(
        mem_2__0_), .QN(n635) );
  FD1S mem_reg_1__35_ ( .D(n445), .TI(mem_1__34_), .TE(test_se), .CP(n23), .Q(
        mem_1__35_), .QN(n670) );
  FD1S mem_reg_1__34_ ( .D(n444), .TI(mem_1__33_), .TE(test_se), .CP(n23), .Q(
        mem_1__34_), .QN(n669) );
  FD1S mem_reg_1__33_ ( .D(n443), .TI(mem_1__32_), .TE(test_se), .CP(n23), .Q(
        mem_1__33_), .QN(n668) );
  FD1S mem_reg_1__32_ ( .D(n442), .TI(mem_1__31_), .TE(test_se), .CP(n23), .Q(
        mem_1__32_), .QN(n667) );
  FD1S mem_reg_1__31_ ( .D(n441), .TI(mem_1__30_), .TE(test_se), .CP(n23), .Q(
        mem_1__31_), .QN(n666) );
  FD1S mem_reg_1__30_ ( .D(n440), .TI(mem_1__29_), .TE(test_se), .CP(n22), .Q(
        mem_1__30_), .QN(n665) );
  FD1S mem_reg_1__29_ ( .D(n439), .TI(mem_1__28_), .TE(test_se), .CP(n22), .Q(
        mem_1__29_), .QN(n664) );
  FD1S mem_reg_1__28_ ( .D(n438), .TI(mem_1__27_), .TE(test_se), .CP(n22), .Q(
        mem_1__28_), .QN(n663) );
  FD1S mem_reg_1__27_ ( .D(n437), .TI(mem_1__26_), .TE(test_se), .CP(n22), .Q(
        mem_1__27_), .QN(n662) );
  FD1S mem_reg_1__26_ ( .D(n436), .TI(mem_1__25_), .TE(test_se), .CP(n22), .Q(
        mem_1__26_), .QN(n661) );
  FD1S mem_reg_1__25_ ( .D(n435), .TI(mem_1__24_), .TE(test_se), .CP(n22), .Q(
        mem_1__25_), .QN(n660) );
  FD1S mem_reg_1__24_ ( .D(n434), .TI(mem_1__23_), .TE(test_se), .CP(n22), .Q(
        mem_1__24_), .QN(n659) );
  FD1S mem_reg_1__23_ ( .D(n433), .TI(mem_1__22_), .TE(test_se), .CP(n22), .Q(
        mem_1__23_), .QN(n658) );
  FD1S mem_reg_1__22_ ( .D(n432), .TI(mem_1__21_), .TE(test_se), .CP(n22), .Q(
        mem_1__22_), .QN(n657) );
  FD1S mem_reg_1__21_ ( .D(n431), .TI(mem_1__20_), .TE(test_se), .CP(n22), .Q(
        mem_1__21_), .QN(n656) );
  FD1S mem_reg_1__20_ ( .D(n430), .TI(mem_1__19_), .TE(test_se), .CP(n22), .Q(
        mem_1__20_), .QN(n655) );
  FD1S mem_reg_1__19_ ( .D(n429), .TI(mem_1__18_), .TE(test_se), .CP(n22), .Q(
        mem_1__19_), .QN(n654) );
  FD1S mem_reg_1__18_ ( .D(n428), .TI(mem_1__17_), .TE(test_se), .CP(n21), .Q(
        mem_1__18_), .QN(n653) );
  FD1S mem_reg_1__17_ ( .D(n427), .TI(mem_1__16_), .TE(test_se), .CP(n21), .Q(
        mem_1__17_), .QN(n652) );
  FD1S mem_reg_1__16_ ( .D(n426), .TI(mem_1__15_), .TE(test_se), .CP(n21), .Q(
        mem_1__16_), .QN(n651) );
  FD1S mem_reg_1__15_ ( .D(n425), .TI(mem_1__14_), .TE(test_se), .CP(n21), .Q(
        mem_1__15_), .QN(n650) );
  FD1S mem_reg_1__14_ ( .D(n424), .TI(mem_1__13_), .TE(test_se), .CP(n21), .Q(
        mem_1__14_), .QN(n649) );
  FD1S mem_reg_1__13_ ( .D(n423), .TI(mem_1__12_), .TE(test_se), .CP(n21), .Q(
        mem_1__13_), .QN(n648) );
  FD1S mem_reg_1__12_ ( .D(n422), .TI(mem_1__11_), .TE(test_se), .CP(n21), .Q(
        mem_1__12_), .QN(n647) );
  FD1S mem_reg_1__11_ ( .D(n421), .TI(mem_1__10_), .TE(test_se), .CP(n21), .Q(
        mem_1__11_), .QN(n646) );
  FD1S mem_reg_1__10_ ( .D(n420), .TI(mem_1__9_), .TE(test_se), .CP(n21), .Q(
        mem_1__10_), .QN(n645) );
  FD1S mem_reg_1__9_ ( .D(n419), .TI(mem_1__8_), .TE(test_se), .CP(n21), .Q(
        mem_1__9_), .QN(n644) );
  FD1S mem_reg_1__8_ ( .D(n418), .TI(mem_1__7_), .TE(test_se), .CP(n21), .Q(
        mem_1__8_), .QN(n643) );
  FD1S mem_reg_1__7_ ( .D(n417), .TI(test_si2), .TE(test_se), .CP(n21), .Q(
        mem_1__7_), .QN(n642) );
  FD1S mem_reg_1__6_ ( .D(n416), .TI(mem_1__5_), .TE(test_se), .CP(n20), .Q(
        test_so1), .QN(n641) );
  FD1S mem_reg_1__5_ ( .D(n415), .TI(mem_1__4_), .TE(test_se), .CP(n20), .Q(
        mem_1__5_), .QN(n640) );
  FD1S mem_reg_1__4_ ( .D(n414), .TI(mem_1__3_), .TE(test_se), .CP(n20), .Q(
        mem_1__4_), .QN(n639) );
  FD1S mem_reg_1__3_ ( .D(n413), .TI(mem_1__2_), .TE(test_se), .CP(n20), .Q(
        mem_1__3_), .QN(n638) );
  FD1S mem_reg_1__2_ ( .D(n412), .TI(mem_1__1_), .TE(test_se), .CP(n20), .Q(
        mem_1__2_), .QN(n637) );
  FD1S mem_reg_1__1_ ( .D(n411), .TI(mem_1__0_), .TE(test_se), .CP(n20), .Q(
        mem_1__1_), .QN(n636) );
  FD1S mem_reg_1__0_ ( .D(n446), .TI(mem_0__35_), .TE(test_se), .CP(n23), .Q(
        mem_1__0_), .QN(n671) );
  FD1S mem_reg_0__35_ ( .D(n481), .TI(mem_0__34_), .TE(test_se), .CP(n26), .Q(
        mem_0__35_), .QN(n706) );
  FD1S mem_reg_0__34_ ( .D(n480), .TI(mem_0__33_), .TE(test_se), .CP(n26), .Q(
        mem_0__34_), .QN(n705) );
  FD1S mem_reg_0__33_ ( .D(n479), .TI(mem_0__32_), .TE(test_se), .CP(n26), .Q(
        mem_0__33_), .QN(n704) );
  FD1S mem_reg_0__32_ ( .D(n478), .TI(mem_0__31_), .TE(test_se), .CP(n26), .Q(
        mem_0__32_), .QN(n703) );
  FD1S mem_reg_0__31_ ( .D(n477), .TI(mem_0__30_), .TE(test_se), .CP(n26), .Q(
        mem_0__31_), .QN(n702) );
  FD1S mem_reg_0__30_ ( .D(n476), .TI(mem_0__29_), .TE(test_se), .CP(n25), .Q(
        mem_0__30_), .QN(n701) );
  FD1S mem_reg_0__29_ ( .D(n475), .TI(mem_0__28_), .TE(test_se), .CP(n25), .Q(
        mem_0__29_), .QN(n700) );
  FD1S mem_reg_0__28_ ( .D(n474), .TI(mem_0__27_), .TE(test_se), .CP(n25), .Q(
        mem_0__28_), .QN(n699) );
  FD1S mem_reg_0__27_ ( .D(n473), .TI(mem_0__26_), .TE(test_se), .CP(n25), .Q(
        mem_0__27_), .QN(n698) );
  FD1S mem_reg_0__26_ ( .D(n472), .TI(mem_0__25_), .TE(test_se), .CP(n25), .Q(
        mem_0__26_), .QN(n697) );
  FD1S mem_reg_0__25_ ( .D(n471), .TI(mem_0__24_), .TE(test_se), .CP(n25), .Q(
        mem_0__25_), .QN(n696) );
  FD1S mem_reg_0__24_ ( .D(n470), .TI(mem_0__23_), .TE(test_se), .CP(n25), .Q(
        mem_0__24_), .QN(n695) );
  FD1S mem_reg_0__23_ ( .D(n469), .TI(mem_0__22_), .TE(test_se), .CP(n25), .Q(
        mem_0__23_), .QN(n694) );
  FD1S mem_reg_0__22_ ( .D(n468), .TI(mem_0__21_), .TE(test_se), .CP(n25), .Q(
        mem_0__22_), .QN(n693) );
  FD1S mem_reg_0__21_ ( .D(n467), .TI(mem_0__20_), .TE(test_se), .CP(n25), .Q(
        mem_0__21_), .QN(n692) );
  FD1S mem_reg_0__20_ ( .D(n466), .TI(mem_0__19_), .TE(test_se), .CP(n25), .Q(
        mem_0__20_), .QN(n691) );
  FD1S mem_reg_0__19_ ( .D(n465), .TI(mem_0__18_), .TE(test_se), .CP(n25), .Q(
        mem_0__19_), .QN(n690) );
  FD1S mem_reg_0__18_ ( .D(n464), .TI(mem_0__17_), .TE(test_se), .CP(n24), .Q(
        mem_0__18_), .QN(n689) );
  FD1S mem_reg_0__17_ ( .D(n463), .TI(mem_0__16_), .TE(test_se), .CP(n24), .Q(
        mem_0__17_), .QN(n688) );
  FD1S mem_reg_0__16_ ( .D(n462), .TI(mem_0__15_), .TE(test_se), .CP(n24), .Q(
        mem_0__16_), .QN(n687) );
  FD1S mem_reg_0__15_ ( .D(n461), .TI(mem_0__14_), .TE(test_se), .CP(n24), .Q(
        mem_0__15_), .QN(n686) );
  FD1S mem_reg_0__14_ ( .D(n460), .TI(mem_0__13_), .TE(test_se), .CP(n24), .Q(
        mem_0__14_), .QN(n685) );
  FD1S mem_reg_0__13_ ( .D(n459), .TI(mem_0__12_), .TE(test_se), .CP(n24), .Q(
        mem_0__13_), .QN(n684) );
  FD1S mem_reg_0__12_ ( .D(n458), .TI(mem_0__11_), .TE(test_se), .CP(n24), .Q(
        mem_0__12_), .QN(n683) );
  FD1S mem_reg_0__11_ ( .D(n457), .TI(mem_0__10_), .TE(test_se), .CP(n24), .Q(
        mem_0__11_), .QN(n682) );
  FD1S mem_reg_0__10_ ( .D(n456), .TI(mem_0__9_), .TE(test_se), .CP(n24), .Q(
        mem_0__10_), .QN(n681) );
  FD1S mem_reg_0__9_ ( .D(n455), .TI(mem_0__8_), .TE(test_se), .CP(n24), .Q(
        mem_0__9_), .QN(n680) );
  FD1S mem_reg_0__8_ ( .D(n454), .TI(mem_0__7_), .TE(test_se), .CP(n24), .Q(
        mem_0__8_), .QN(n679) );
  FD1S mem_reg_0__7_ ( .D(n453), .TI(mem_0__6_), .TE(test_se), .CP(n24), .Q(
        mem_0__7_), .QN(n678) );
  FD1S mem_reg_0__6_ ( .D(n452), .TI(mem_0__5_), .TE(test_se), .CP(n23), .Q(
        mem_0__6_), .QN(n677) );
  FD1S mem_reg_0__5_ ( .D(n451), .TI(mem_0__4_), .TE(test_se), .CP(n23), .Q(
        mem_0__5_), .QN(n676) );
  FD1S mem_reg_0__4_ ( .D(n450), .TI(mem_0__3_), .TE(test_se), .CP(n23), .Q(
        mem_0__4_), .QN(n675) );
  FD1S mem_reg_0__3_ ( .D(n449), .TI(mem_0__2_), .TE(test_se), .CP(n23), .Q(
        mem_0__3_), .QN(n674) );
  FD1S mem_reg_0__2_ ( .D(n448), .TI(mem_0__1_), .TE(test_se), .CP(n23), .Q(
        mem_0__2_), .QN(n673) );
  FD1S mem_reg_0__1_ ( .D(n447), .TI(mem_0__0_), .TE(test_se), .CP(n23), .Q(
        mem_0__1_), .QN(n672) );
  FD1S mem_reg_0__0_ ( .D(n482), .TI(grey_wr_ptr[2]), .TE(test_se), .CP(n26), 
        .Q(mem_0__0_), .QN(n707) );
  FD1S rd_data_q_reg_35_ ( .D(rd_data_c[35]), .TI(rd_data[34]), .TE(test_se), 
        .CP(n8), .Q(rd_data[35]) );
  FD1S rd_data_q_reg_28_ ( .D(rd_data_c[28]), .TI(rd_data[27]), .TE(test_se), 
        .CP(n8), .Q(rd_data[28]) );
  FD1S rd_data_q_reg_25_ ( .D(rd_data_c[25]), .TI(rd_data[24]), .TE(test_se), 
        .CP(n7), .Q(rd_data[25]) );
  FD1S rd_data_q_reg_6_ ( .D(rd_data_c[6]), .TI(rd_data[5]), .TE(test_se), 
        .CP(n6), .Q(rd_data[6]) );
  FD4S empty_q_reg ( .D(n333), .TI(test_si5), .TE(test_se), .CP(n9), .SD(
        rd_reset_n), .Q(empty), .QN(n561) );
  FD2S grey_wr_ptr_reg_2_ ( .D(n337), .TI(grey_wr_ptr[1]), .TE(test_se), .CP(
        n14), .CD(wr_reset_n), .Q(grey_wr_ptr[2]), .QN(n563) );
  FD2S grey_rd_ptr_reg_2_ ( .D(n486), .TI(grey_rd_ptr_dly[1]), .TE(test_se), 
        .CP(n8), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[2]), .QN(n709) );
  FD2S grey_rd_ptr_reg_1_ ( .D(n484), .TI(grey_rd_ptr_dly[0]), .TE(test_se), 
        .CP(n8), .CD(rd_reset_n), .Q(grey_rd_ptr_dly[1]), .QN(n708) );
  FD1S rd_data_q_reg_34_ ( .D(rd_data_c[34]), .TI(rd_data[33]), .TE(test_se), 
        .CP(n8), .Q(rd_data[34]) );
  FD1S rd_data_q_reg_30_ ( .D(rd_data_c[30]), .TI(rd_data[29]), .TE(test_se), 
        .CP(n8), .Q(rd_data[30]) );
  FD1S rd_data_q_reg_29_ ( .D(rd_data_c[29]), .TI(rd_data[28]), .TE(test_se), 
        .CP(n8), .Q(rd_data[29]) );
  FD1S rd_data_q_reg_26_ ( .D(rd_data_c[26]), .TI(rd_data[25]), .TE(test_se), 
        .CP(n7), .Q(rd_data[26]) );
  FD1S rd_data_q_reg_24_ ( .D(rd_data_c[24]), .TI(rd_data[23]), .TE(test_se), 
        .CP(n7), .Q(rd_data[24]) );
  FD1S rd_data_q_reg_3_ ( .D(rd_data_c[3]), .TI(rd_data[2]), .TE(test_se), 
        .CP(n5), .Q(rd_data[3]) );
  FD1S rd_data_q_reg_2_ ( .D(rd_data_c[2]), .TI(rd_data[1]), .TE(test_se), 
        .CP(n5), .Q(rd_data[2]) );
  FD2S grey_wr_ptr_reg_1_ ( .D(n335), .TI(grey_wr_ptr[0]), .TE(test_se), .CP(
        n14), .CD(wr_reset_n), .Q(grey_wr_ptr[1]) );
  FD2S rd_ptr_reg_2_ ( .D(n487), .TI(N46), .TE(test_se), .CP(n8), .CD(
        rd_reset_n), .Q(n712), .QN(n3) );
  FD2S sync_rd_ptr_1_reg_1_ ( .D(sync_rd_ptr_0[1]), .TI(sync_rd_ptr_1[0]), 
        .TE(test_se), .CP(n26), .CD(wr_reset_n), .Q(sync_rd_ptr_1[1]), .QN(
        n711) );
  FD2S sync_rd_ptr_1_reg_0_ ( .D(sync_rd_ptr_0[0]), .TI(sync_rd_ptr_0[2]), 
        .TE(test_se), .CP(n26), .CD(wr_reset_n), .Q(sync_rd_ptr_1[0]) );
  FD2S full_q_reg ( .D(n334), .TI(test_si1), .TE(test_se), .CP(n27), .CD(
        wr_reset_n), .Q(full), .QN(n562) );
  FD2S sync_wr_ptr_1_reg_0_ ( .D(sync_wr_ptr_0[0]), .TI(sync_wr_ptr_0[2]), 
        .TE(test_se), .CP(n5), .CD(rd_reset_n), .Q(sync_wr_ptr_1_0_) );
  FD1S rd_data_q_reg_33_ ( .D(rd_data_c[33]), .TI(rd_data[32]), .TE(test_se), 
        .CP(n8), .Q(rd_data[33]) );
  FD1S rd_data_q_reg_32_ ( .D(rd_data_c[32]), .TI(rd_data[31]), .TE(test_se), 
        .CP(n8), .Q(rd_data[32]) );
  FD1S rd_data_q_reg_31_ ( .D(rd_data_c[31]), .TI(rd_data[30]), .TE(test_se), 
        .CP(n8), .Q(rd_data[31]) );
  FD1S rd_data_q_reg_23_ ( .D(rd_data_c[23]), .TI(rd_data[22]), .TE(test_se), 
        .CP(n7), .Q(rd_data[23]) );
  FD1S rd_data_q_reg_22_ ( .D(rd_data_c[22]), .TI(rd_data[21]), .TE(test_se), 
        .CP(n7), .Q(rd_data[22]) );
  FD1S rd_data_q_reg_21_ ( .D(rd_data_c[21]), .TI(rd_data[20]), .TE(test_se), 
        .CP(n7), .Q(rd_data[21]) );
  FD1S rd_data_q_reg_20_ ( .D(rd_data_c[20]), .TI(rd_data[19]), .TE(test_se), 
        .CP(n7), .Q(rd_data[20]) );
  FD1S rd_data_q_reg_19_ ( .D(rd_data_c[19]), .TI(rd_data[18]), .TE(test_se), 
        .CP(n7), .Q(rd_data[19]) );
  FD1S rd_data_q_reg_18_ ( .D(rd_data_c[18]), .TI(rd_data[17]), .TE(test_se), 
        .CP(n7), .Q(rd_data[18]) );
  FD1S rd_data_q_reg_17_ ( .D(rd_data_c[17]), .TI(rd_data[16]), .TE(test_se), 
        .CP(n7), .Q(rd_data[17]) );
  FD1S rd_data_q_reg_16_ ( .D(rd_data_c[16]), .TI(rd_data[15]), .TE(test_se), 
        .CP(n7), .Q(rd_data[16]) );
  FD1S rd_data_q_reg_15_ ( .D(rd_data_c[15]), .TI(rd_data[14]), .TE(test_se), 
        .CP(n6), .Q(rd_data[15]) );
  FD1S rd_data_q_reg_14_ ( .D(rd_data_c[14]), .TI(rd_data[13]), .TE(test_se), 
        .CP(n6), .Q(rd_data[14]) );
  FD1S rd_data_q_reg_13_ ( .D(rd_data_c[13]), .TI(test_si6), .TE(test_se), 
        .CP(n6), .Q(rd_data[13]) );
  FD1S rd_data_q_reg_12_ ( .D(rd_data_c[12]), .TI(rd_data[11]), .TE(test_se), 
        .CP(n6), .Q(rd_data[12]) );
  FD1S rd_data_q_reg_11_ ( .D(rd_data_c[11]), .TI(rd_data[10]), .TE(test_se), 
        .CP(n6), .Q(rd_data[11]) );
  FD1S rd_data_q_reg_7_ ( .D(rd_data_c[7]), .TI(rd_data[6]), .TE(test_se), 
        .CP(n6), .Q(rd_data[7]) );
  FD1S rd_data_q_reg_5_ ( .D(rd_data_c[5]), .TI(rd_data[4]), .TE(test_se), 
        .CP(n6), .Q(rd_data[5]) );
  FD1S rd_data_q_reg_4_ ( .D(rd_data_c[4]), .TI(rd_data[3]), .TE(test_se), 
        .CP(n6), .Q(rd_data[4]) );
  FD1S rd_data_q_reg_1_ ( .D(rd_data_c[1]), .TI(rd_data[0]), .TE(test_se), 
        .CP(n5), .Q(rd_data[1]) );
  FD1S rd_data_q_reg_0_ ( .D(rd_data_c[0]), .TI(grey_rd_ptr_dly[2]), .TE(
        test_se), .CP(n5), .Q(rd_data[0]) );
  FD2S wr_ptr_reg_2_ ( .D(n338), .TI(wr_ptr[1]), .TE(test_se), .CP(n14), .CD(
        wr_reset_n), .Q(test_so4), .QN(n2) );
  FD2S grey_wr_ptr_reg_0_ ( .D(n336), .TI(full), .TE(test_se), .CP(n14), .CD(
        wr_reset_n), .Q(grey_wr_ptr[0]) );
  FD2S grey_rd_ptr_reg_0_ ( .D(n485), .TI(empty), .TE(test_se), .CP(n8), .CD(
        rd_reset_n), .Q(grey_rd_ptr_dly[0]) );
  FD1S rd_data_q_reg_27_ ( .D(rd_data_c[27]), .TI(rd_data[26]), .TE(test_se), 
        .CP(n7), .Q(rd_data[27]) );
  FD1S rd_data_q_reg_10_ ( .D(rd_data_c[10]), .TI(rd_data[9]), .TE(test_se), 
        .CP(n6), .Q(rd_data[10]) );
  FD1S rd_data_q_reg_9_ ( .D(rd_data_c[9]), .TI(rd_data[8]), .TE(test_se), 
        .CP(n6), .Q(rd_data[9]) );
  FD1S rd_data_q_reg_8_ ( .D(rd_data_c[8]), .TI(rd_data[7]), .TE(test_se), 
        .CP(n6), .Q(rd_data[8]) );
  FD2S sync_rd_ptr_1_reg_2_ ( .D(sync_rd_ptr_0[2]), .TI(sync_rd_ptr_1[1]), 
        .TE(test_se), .CP(n26), .CD(wr_reset_n), .Q(sync_rd_ptr_1[2]) );
  FD2S sync_wr_ptr_1_reg_2_ ( .D(sync_wr_ptr_0[2]), .TI(n716), .TE(test_se), 
        .CP(n5), .CD(rd_reset_n), .Q(test_so5) );
  FD2S wr_ptr_reg_1_ ( .D(n483), .TI(wr_ptr[0]), .TE(test_se), .CP(n14), .CD(
        wr_reset_n), .Q(wr_ptr[1]), .QN(n1) );
  FD2S rd_ptr_reg_0_ ( .D(n489), .TI(rd_data[35]), .TE(test_se), .CP(n5), .CD(
        rd_reset_n), .Q(N45), .QN(n248) );
  FD2S rd_ptr_reg_1_ ( .D(n488), .TI(N45), .TE(test_se), .CP(n5), .CD(
        rd_reset_n), .Q(N46), .QN(n246) );
  FD2S wr_ptr_reg_0_ ( .D(n714), .TI(sync_rd_ptr_1[2]), .TE(test_se), .CP(n14), 
        .CD(wr_reset_n), .Q(wr_ptr[0]), .QN(n4) );
  FD2S sync_rd_ptr_0_reg_2_ ( .D(grey_rd_ptr_dly[2]), .TI(sync_rd_ptr_0[1]), 
        .TE(test_se), .CP(n26), .CD(wr_reset_n), .Q(sync_rd_ptr_0[2]) );
  FD2S sync_rd_ptr_0_reg_1_ ( .D(grey_rd_ptr_dly[1]), .TI(sync_rd_ptr_0[0]), 
        .TE(test_se), .CP(n26), .CD(wr_reset_n), .Q(sync_rd_ptr_0[1]) );
  FD2S sync_rd_ptr_0_reg_0_ ( .D(grey_rd_ptr_dly[0]), .TI(mem_3__35_), .TE(
        test_se), .CP(n26), .CD(wr_reset_n), .Q(sync_rd_ptr_0[0]) );
  FD2S sync_wr_ptr_0_reg_2_ ( .D(grey_wr_ptr[2]), .TI(sync_wr_ptr_0[1]), .TE(
        test_se), .CP(n5), .CD(rd_reset_n), .Q(sync_wr_ptr_0[2]) );
  FD2S sync_wr_ptr_0_reg_1_ ( .D(grey_wr_ptr[1]), .TI(sync_wr_ptr_0[0]), .TE(
        test_se), .CP(n5), .CD(rd_reset_n), .Q(sync_wr_ptr_0[1]) );
  FD2S sync_wr_ptr_0_reg_0_ ( .D(grey_wr_ptr[0]), .TI(n712), .TE(test_se), 
        .CP(n5), .CD(rd_reset_n), .Q(sync_wr_ptr_0[0]) );
  IVP U209 ( .A(n29), .Z(n24) );
  IVP U210 ( .A(n28), .Z(n25) );
  IVP U211 ( .A(n28), .Z(n26) );
  IVP U212 ( .A(n30), .Z(n21) );
  IVP U213 ( .A(n29), .Z(n22) );
  IVP U214 ( .A(n29), .Z(n23) );
  IVP U215 ( .A(n237), .Z(n18) );
  IVP U216 ( .A(n30), .Z(n19) );
  IVP U217 ( .A(n30), .Z(n20) );
  IVP U218 ( .A(n238), .Z(n15) );
  IVP U219 ( .A(n237), .Z(n16) );
  IVP U220 ( .A(n237), .Z(n17) );
  IVP U221 ( .A(n238), .Z(n14) );
  IVP U222 ( .A(n28), .Z(n27) );
  IVP U223 ( .A(n240), .Z(n28) );
  IVP U224 ( .A(n240), .Z(n29) );
  IVP U225 ( .A(n239), .Z(n30) );
  IVP U226 ( .A(n239), .Z(n237) );
  IVP U227 ( .A(n239), .Z(n238) );
  IVP U228 ( .A(n11), .Z(n6) );
  IVP U229 ( .A(n10), .Z(n7) );
  IVP U230 ( .A(n10), .Z(n8) );
  IVP U231 ( .A(n11), .Z(n5) );
  IVP U232 ( .A(n10), .Z(n9) );
  IVP U233 ( .A(n241), .Z(n239) );
  IVP U234 ( .A(n12), .Z(n10) );
  IVP U235 ( .A(n241), .Z(n240) );
  IVP U236 ( .A(n12), .Z(n11) );
  IVP U237 ( .A(wr_clk), .Z(n241) );
  IVP U238 ( .A(n13), .Z(n12) );
  IVP U239 ( .A(rd_clk), .Z(n13) );
  NR2 U240 ( .A(n246), .B(N45), .Z(n315) );
  NR2 U241 ( .A(n246), .B(n248), .Z(n314) );
  AO2 U242 ( .A(mem_2__0_), .B(n315), .C(mem_3__0_), .D(n314), .Z(n243) );
  NR2 U243 ( .A(N45), .B(N46), .Z(n317) );
  NR2 U244 ( .A(n248), .B(N46), .Z(n316) );
  AO2 U245 ( .A(mem_0__0_), .B(n317), .C(mem_1__0_), .D(n316), .Z(n242) );
  ND2 U246 ( .A(n243), .B(n242), .Z(rd_data_c[0]) );
  AO2 U247 ( .A(mem_2__1_), .B(n315), .C(mem_3__1_), .D(n314), .Z(n245) );
  AO2 U248 ( .A(mem_0__1_), .B(n317), .C(mem_1__1_), .D(n316), .Z(n244) );
  ND2 U249 ( .A(n245), .B(n244), .Z(rd_data_c[1]) );
  AO2 U250 ( .A(mem_2__2_), .B(n315), .C(mem_3__2_), .D(n314), .Z(n249) );
  AO2 U251 ( .A(mem_0__2_), .B(n317), .C(mem_1__2_), .D(n316), .Z(n247) );
  ND2 U252 ( .A(n249), .B(n247), .Z(rd_data_c[2]) );
  AO2 U253 ( .A(mem_2__3_), .B(n315), .C(mem_3__3_), .D(n314), .Z(n251) );
  AO2 U254 ( .A(mem_0__3_), .B(n317), .C(mem_1__3_), .D(n316), .Z(n250) );
  ND2 U255 ( .A(n251), .B(n250), .Z(rd_data_c[3]) );
  AO2 U256 ( .A(mem_2__4_), .B(n315), .C(mem_3__4_), .D(n314), .Z(n253) );
  AO2 U257 ( .A(mem_0__4_), .B(n317), .C(mem_1__4_), .D(n316), .Z(n252) );
  ND2 U258 ( .A(n253), .B(n252), .Z(rd_data_c[4]) );
  AO2 U259 ( .A(mem_2__5_), .B(n315), .C(mem_3__5_), .D(n314), .Z(n255) );
  AO2 U260 ( .A(mem_0__5_), .B(n317), .C(mem_1__5_), .D(n316), .Z(n254) );
  ND2 U261 ( .A(n255), .B(n254), .Z(rd_data_c[5]) );
  AO2 U262 ( .A(mem_2__6_), .B(n315), .C(mem_3__6_), .D(n314), .Z(n257) );
  AO2 U263 ( .A(mem_0__6_), .B(n317), .C(test_so1), .D(n316), .Z(n256) );
  ND2 U264 ( .A(n257), .B(n256), .Z(rd_data_c[6]) );
  AO2 U265 ( .A(mem_2__7_), .B(n315), .C(mem_3__7_), .D(n314), .Z(n259) );
  AO2 U266 ( .A(mem_0__7_), .B(n317), .C(mem_1__7_), .D(n316), .Z(n258) );
  ND2 U267 ( .A(n259), .B(n258), .Z(rd_data_c[7]) );
  AO2 U268 ( .A(mem_2__8_), .B(n315), .C(mem_3__8_), .D(n314), .Z(n261) );
  AO2 U269 ( .A(mem_0__8_), .B(n317), .C(mem_1__8_), .D(n316), .Z(n260) );
  ND2 U270 ( .A(n261), .B(n260), .Z(rd_data_c[8]) );
  AO2 U271 ( .A(mem_2__9_), .B(n315), .C(mem_3__9_), .D(n314), .Z(n263) );
  AO2 U272 ( .A(mem_0__9_), .B(n317), .C(mem_1__9_), .D(n316), .Z(n262) );
  ND2 U273 ( .A(n263), .B(n262), .Z(rd_data_c[9]) );
  AO2 U274 ( .A(mem_2__10_), .B(n315), .C(mem_3__10_), .D(n314), .Z(n265) );
  AO2 U275 ( .A(mem_0__10_), .B(n317), .C(mem_1__10_), .D(n316), .Z(n264) );
  ND2 U276 ( .A(n265), .B(n264), .Z(rd_data_c[10]) );
  AO2 U277 ( .A(mem_2__11_), .B(n315), .C(mem_3__11_), .D(n314), .Z(n267) );
  AO2 U278 ( .A(mem_0__11_), .B(n317), .C(mem_1__11_), .D(n316), .Z(n266) );
  ND2 U279 ( .A(n267), .B(n266), .Z(rd_data_c[11]) );
  AO2 U280 ( .A(mem_2__12_), .B(n315), .C(mem_3__12_), .D(n314), .Z(n269) );
  AO2 U281 ( .A(mem_0__12_), .B(n317), .C(mem_1__12_), .D(n316), .Z(n268) );
  ND2 U282 ( .A(n269), .B(n268), .Z(rd_data_c[12]) );
  AO2 U283 ( .A(mem_2__13_), .B(n315), .C(mem_3__13_), .D(n314), .Z(n271) );
  AO2 U284 ( .A(mem_0__13_), .B(n317), .C(mem_1__13_), .D(n316), .Z(n270) );
  ND2 U285 ( .A(n271), .B(n270), .Z(rd_data_c[13]) );
  AO2 U286 ( .A(mem_2__14_), .B(n315), .C(mem_3__14_), .D(n314), .Z(n273) );
  AO2 U287 ( .A(mem_0__14_), .B(n317), .C(mem_1__14_), .D(n316), .Z(n272) );
  ND2 U288 ( .A(n273), .B(n272), .Z(rd_data_c[14]) );
  AO2 U289 ( .A(mem_2__15_), .B(n315), .C(mem_3__15_), .D(n314), .Z(n275) );
  AO2 U290 ( .A(mem_0__15_), .B(n317), .C(mem_1__15_), .D(n316), .Z(n274) );
  ND2 U291 ( .A(n275), .B(n274), .Z(rd_data_c[15]) );
  AO2 U292 ( .A(mem_2__16_), .B(n315), .C(mem_3__16_), .D(n314), .Z(n277) );
  AO2 U293 ( .A(mem_0__16_), .B(n317), .C(mem_1__16_), .D(n316), .Z(n276) );
  ND2 U294 ( .A(n277), .B(n276), .Z(rd_data_c[16]) );
  AO2 U295 ( .A(mem_2__17_), .B(n315), .C(mem_3__17_), .D(n314), .Z(n279) );
  AO2 U296 ( .A(mem_0__17_), .B(n317), .C(mem_1__17_), .D(n316), .Z(n278) );
  ND2 U297 ( .A(n279), .B(n278), .Z(rd_data_c[17]) );
  AO2 U298 ( .A(test_so2), .B(n315), .C(mem_3__18_), .D(n314), .Z(n281) );
  AO2 U299 ( .A(mem_0__18_), .B(n317), .C(mem_1__18_), .D(n316), .Z(n280) );
  ND2 U300 ( .A(n281), .B(n280), .Z(rd_data_c[18]) );
  AO2 U301 ( .A(mem_2__19_), .B(n315), .C(mem_3__19_), .D(n314), .Z(n283) );
  AO2 U302 ( .A(mem_0__19_), .B(n317), .C(mem_1__19_), .D(n316), .Z(n282) );
  ND2 U303 ( .A(n283), .B(n282), .Z(rd_data_c[19]) );
  AO2 U304 ( .A(mem_2__20_), .B(n315), .C(mem_3__20_), .D(n314), .Z(n285) );
  AO2 U305 ( .A(mem_0__20_), .B(n317), .C(mem_1__20_), .D(n316), .Z(n284) );
  ND2 U306 ( .A(n285), .B(n284), .Z(rd_data_c[20]) );
  AO2 U307 ( .A(mem_2__21_), .B(n315), .C(mem_3__21_), .D(n314), .Z(n287) );
  AO2 U308 ( .A(mem_0__21_), .B(n317), .C(mem_1__21_), .D(n316), .Z(n286) );
  ND2 U309 ( .A(n287), .B(n286), .Z(rd_data_c[21]) );
  AO2 U310 ( .A(mem_2__22_), .B(n315), .C(mem_3__22_), .D(n314), .Z(n289) );
  AO2 U311 ( .A(mem_0__22_), .B(n317), .C(mem_1__22_), .D(n316), .Z(n288) );
  ND2 U312 ( .A(n289), .B(n288), .Z(rd_data_c[22]) );
  AO2 U313 ( .A(mem_2__23_), .B(n315), .C(mem_3__23_), .D(n314), .Z(n291) );
  AO2 U314 ( .A(mem_0__23_), .B(n317), .C(mem_1__23_), .D(n316), .Z(n290) );
  ND2 U315 ( .A(n291), .B(n290), .Z(rd_data_c[23]) );
  AO2 U316 ( .A(mem_2__24_), .B(n315), .C(mem_3__24_), .D(n314), .Z(n293) );
  AO2 U317 ( .A(mem_0__24_), .B(n317), .C(mem_1__24_), .D(n316), .Z(n292) );
  ND2 U318 ( .A(n293), .B(n292), .Z(rd_data_c[24]) );
  AO2 U319 ( .A(mem_2__25_), .B(n315), .C(mem_3__25_), .D(n314), .Z(n295) );
  AO2 U320 ( .A(mem_0__25_), .B(n317), .C(mem_1__25_), .D(n316), .Z(n294) );
  ND2 U321 ( .A(n295), .B(n294), .Z(rd_data_c[25]) );
  AO2 U322 ( .A(mem_2__26_), .B(n315), .C(mem_3__26_), .D(n314), .Z(n297) );
  AO2 U323 ( .A(mem_0__26_), .B(n317), .C(mem_1__26_), .D(n316), .Z(n296) );
  ND2 U324 ( .A(n297), .B(n296), .Z(rd_data_c[26]) );
  AO2 U325 ( .A(mem_2__27_), .B(n315), .C(mem_3__27_), .D(n314), .Z(n299) );
  AO2 U326 ( .A(mem_0__27_), .B(n317), .C(mem_1__27_), .D(n316), .Z(n298) );
  ND2 U327 ( .A(n299), .B(n298), .Z(rd_data_c[27]) );
  AO2 U328 ( .A(mem_2__28_), .B(n315), .C(mem_3__28_), .D(n314), .Z(n301) );
  AO2 U329 ( .A(mem_0__28_), .B(n317), .C(mem_1__28_), .D(n316), .Z(n300) );
  ND2 U330 ( .A(n301), .B(n300), .Z(rd_data_c[28]) );
  AO2 U331 ( .A(mem_2__29_), .B(n315), .C(mem_3__29_), .D(n314), .Z(n303) );
  AO2 U332 ( .A(mem_0__29_), .B(n317), .C(mem_1__29_), .D(n316), .Z(n302) );
  ND2 U333 ( .A(n303), .B(n302), .Z(rd_data_c[29]) );
  AO2 U334 ( .A(mem_2__30_), .B(n315), .C(test_so3), .D(n314), .Z(n305) );
  AO2 U335 ( .A(mem_0__30_), .B(n317), .C(mem_1__30_), .D(n316), .Z(n304) );
  ND2 U336 ( .A(n305), .B(n304), .Z(rd_data_c[30]) );
  AO2 U337 ( .A(mem_2__31_), .B(n315), .C(mem_3__31_), .D(n314), .Z(n307) );
  AO2 U338 ( .A(mem_0__31_), .B(n317), .C(mem_1__31_), .D(n316), .Z(n306) );
  ND2 U339 ( .A(n307), .B(n306), .Z(rd_data_c[31]) );
  AO2 U340 ( .A(mem_2__32_), .B(n315), .C(mem_3__32_), .D(n314), .Z(n309) );
  AO2 U341 ( .A(mem_0__32_), .B(n317), .C(mem_1__32_), .D(n316), .Z(n308) );
  ND2 U342 ( .A(n309), .B(n308), .Z(rd_data_c[32]) );
  AO2 U343 ( .A(mem_2__33_), .B(n315), .C(mem_3__33_), .D(n314), .Z(n311) );
  AO2 U344 ( .A(mem_0__33_), .B(n317), .C(mem_1__33_), .D(n316), .Z(n310) );
  ND2 U345 ( .A(n311), .B(n310), .Z(rd_data_c[33]) );
  AO2 U346 ( .A(mem_2__34_), .B(n315), .C(mem_3__34_), .D(n314), .Z(n313) );
  AO2 U347 ( .A(mem_0__34_), .B(n317), .C(mem_1__34_), .D(n316), .Z(n312) );
  ND2 U348 ( .A(n313), .B(n312), .Z(rd_data_c[34]) );
  AO2 U349 ( .A(mem_2__35_), .B(n315), .C(mem_3__35_), .D(n314), .Z(n319) );
  AO2 U350 ( .A(mem_0__35_), .B(n317), .C(mem_1__35_), .D(n316), .Z(n318) );
  ND2 U351 ( .A(n319), .B(n318), .Z(rd_data_c[35]) );
  EO U352 ( .A(wr_ptr[0]), .B(wr_en), .Z(n714) );
  EO U353 ( .A(N45), .B(rd_en), .Z(n489) );
  AO7 U354 ( .A(rd_en), .B(n246), .C(n320), .Z(n488) );
  AO7 U355 ( .A(rd_en), .B(n3), .C(n321), .Z(n487) );
  AO7 U356 ( .A(rd_en), .B(n709), .C(n321), .Z(n486) );
  AO7 U357 ( .A(n248), .B(n320), .C(n322), .Z(n485) );
  MUX21L U358 ( .A(grey_rd_ptr_dly[0]), .B(n323), .S(rd_en), .Z(n322) );
  NR2 U359 ( .A(n324), .B(N45), .Z(n323) );
  AO7 U360 ( .A(rd_en), .B(n708), .C(n325), .Z(n484) );
  IV U361 ( .A(n326), .Z(n325) );
  AO4 U362 ( .A(n327), .B(n320), .C(n321), .D(n324), .Z(n326) );
  ND2 U363 ( .A(rd_en), .B(n327), .Z(n321) );
  ND2 U364 ( .A(rd_en), .B(n324), .Z(n320) );
  EO U365 ( .A(n246), .B(n248), .Z(n324) );
  EN U366 ( .A(n3), .B(n328), .Z(n327) );
  NR2 U367 ( .A(n246), .B(n248), .Z(n328) );
  AO7 U368 ( .A(wr_en), .B(n1), .C(n329), .Z(n483) );
  MUX21L U369 ( .A(n707), .B(n330), .S(n331), .Z(n482) );
  MUX21L U370 ( .A(n706), .B(n332), .S(n331), .Z(n481) );
  MUX21L U371 ( .A(n705), .B(n490), .S(n331), .Z(n480) );
  MUX21L U372 ( .A(n704), .B(n491), .S(n331), .Z(n479) );
  MUX21L U373 ( .A(n703), .B(n492), .S(n331), .Z(n478) );
  MUX21L U374 ( .A(n702), .B(n493), .S(n331), .Z(n477) );
  MUX21L U375 ( .A(n701), .B(n494), .S(n331), .Z(n476) );
  MUX21L U376 ( .A(n700), .B(n495), .S(n331), .Z(n475) );
  MUX21L U377 ( .A(n699), .B(n496), .S(n331), .Z(n474) );
  MUX21L U378 ( .A(n698), .B(n497), .S(n331), .Z(n473) );
  MUX21L U379 ( .A(n697), .B(n498), .S(n331), .Z(n472) );
  MUX21L U380 ( .A(n696), .B(n499), .S(n331), .Z(n471) );
  MUX21L U381 ( .A(n695), .B(n500), .S(n331), .Z(n470) );
  MUX21L U382 ( .A(n694), .B(n501), .S(n331), .Z(n469) );
  MUX21L U383 ( .A(n693), .B(n502), .S(n331), .Z(n468) );
  MUX21L U384 ( .A(n692), .B(n503), .S(n331), .Z(n467) );
  MUX21L U385 ( .A(n691), .B(n504), .S(n331), .Z(n466) );
  MUX21L U386 ( .A(n690), .B(n505), .S(n331), .Z(n465) );
  MUX21L U387 ( .A(n689), .B(n506), .S(n331), .Z(n464) );
  MUX21L U388 ( .A(n688), .B(n507), .S(n331), .Z(n463) );
  MUX21L U389 ( .A(n687), .B(n508), .S(n331), .Z(n462) );
  MUX21L U390 ( .A(n686), .B(n509), .S(n331), .Z(n461) );
  MUX21L U391 ( .A(n685), .B(n510), .S(n331), .Z(n460) );
  MUX21L U392 ( .A(n684), .B(n511), .S(n331), .Z(n459) );
  MUX21L U393 ( .A(n683), .B(n512), .S(n331), .Z(n458) );
  MUX21L U394 ( .A(n682), .B(n513), .S(n331), .Z(n457) );
  MUX21L U395 ( .A(n681), .B(n514), .S(n331), .Z(n456) );
  MUX21L U396 ( .A(n680), .B(n515), .S(n331), .Z(n455) );
  MUX21L U397 ( .A(n679), .B(n516), .S(n331), .Z(n454) );
  MUX21L U398 ( .A(n678), .B(n517), .S(n331), .Z(n453) );
  MUX21L U399 ( .A(n677), .B(n518), .S(n331), .Z(n452) );
  MUX21L U400 ( .A(n676), .B(n519), .S(n331), .Z(n451) );
  MUX21L U401 ( .A(n675), .B(n520), .S(n331), .Z(n450) );
  MUX21L U402 ( .A(n674), .B(n521), .S(n331), .Z(n449) );
  MUX21L U403 ( .A(n673), .B(n522), .S(n331), .Z(n448) );
  MUX21L U404 ( .A(n672), .B(n523), .S(n331), .Z(n447) );
  NR3 U405 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .C(n524), .Z(n331) );
  MUX21L U406 ( .A(n671), .B(n330), .S(n525), .Z(n446) );
  MUX21L U407 ( .A(n670), .B(n332), .S(n525), .Z(n445) );
  MUX21L U408 ( .A(n669), .B(n490), .S(n525), .Z(n444) );
  MUX21L U409 ( .A(n668), .B(n491), .S(n525), .Z(n443) );
  MUX21L U410 ( .A(n667), .B(n492), .S(n525), .Z(n442) );
  MUX21L U411 ( .A(n666), .B(n493), .S(n525), .Z(n441) );
  MUX21L U412 ( .A(n665), .B(n494), .S(n525), .Z(n440) );
  MUX21L U413 ( .A(n664), .B(n495), .S(n525), .Z(n439) );
  MUX21L U414 ( .A(n663), .B(n496), .S(n525), .Z(n438) );
  MUX21L U415 ( .A(n662), .B(n497), .S(n525), .Z(n437) );
  MUX21L U416 ( .A(n661), .B(n498), .S(n525), .Z(n436) );
  MUX21L U417 ( .A(n660), .B(n499), .S(n525), .Z(n435) );
  MUX21L U418 ( .A(n659), .B(n500), .S(n525), .Z(n434) );
  MUX21L U419 ( .A(n658), .B(n501), .S(n525), .Z(n433) );
  MUX21L U420 ( .A(n657), .B(n502), .S(n525), .Z(n432) );
  MUX21L U421 ( .A(n656), .B(n503), .S(n525), .Z(n431) );
  MUX21L U422 ( .A(n655), .B(n504), .S(n525), .Z(n430) );
  MUX21L U423 ( .A(n654), .B(n505), .S(n525), .Z(n429) );
  MUX21L U424 ( .A(n653), .B(n506), .S(n525), .Z(n428) );
  MUX21L U425 ( .A(n652), .B(n507), .S(n525), .Z(n427) );
  MUX21L U426 ( .A(n651), .B(n508), .S(n525), .Z(n426) );
  MUX21L U427 ( .A(n650), .B(n509), .S(n525), .Z(n425) );
  MUX21L U428 ( .A(n649), .B(n510), .S(n525), .Z(n424) );
  MUX21L U429 ( .A(n648), .B(n511), .S(n525), .Z(n423) );
  MUX21L U430 ( .A(n647), .B(n512), .S(n525), .Z(n422) );
  MUX21L U431 ( .A(n646), .B(n513), .S(n525), .Z(n421) );
  MUX21L U432 ( .A(n645), .B(n514), .S(n525), .Z(n420) );
  MUX21L U433 ( .A(n644), .B(n515), .S(n525), .Z(n419) );
  MUX21L U434 ( .A(n643), .B(n516), .S(n525), .Z(n418) );
  MUX21L U435 ( .A(n642), .B(n517), .S(n525), .Z(n417) );
  MUX21L U436 ( .A(n641), .B(n518), .S(n525), .Z(n416) );
  MUX21L U437 ( .A(n640), .B(n519), .S(n525), .Z(n415) );
  MUX21L U438 ( .A(n639), .B(n520), .S(n525), .Z(n414) );
  MUX21L U439 ( .A(n638), .B(n521), .S(n525), .Z(n413) );
  MUX21L U440 ( .A(n637), .B(n522), .S(n525), .Z(n412) );
  MUX21L U441 ( .A(n636), .B(n523), .S(n525), .Z(n411) );
  NR3 U442 ( .A(n4), .B(wr_ptr[1]), .C(n524), .Z(n525) );
  MUX21L U443 ( .A(n635), .B(n330), .S(n526), .Z(n410) );
  MUX21L U444 ( .A(n634), .B(n332), .S(n526), .Z(n409) );
  MUX21L U445 ( .A(n633), .B(n490), .S(n526), .Z(n408) );
  MUX21L U446 ( .A(n632), .B(n491), .S(n526), .Z(n407) );
  MUX21L U447 ( .A(n631), .B(n492), .S(n526), .Z(n406) );
  MUX21L U448 ( .A(n630), .B(n493), .S(n526), .Z(n405) );
  MUX21L U449 ( .A(n629), .B(n494), .S(n526), .Z(n404) );
  MUX21L U450 ( .A(n628), .B(n495), .S(n526), .Z(n403) );
  MUX21L U451 ( .A(n627), .B(n496), .S(n526), .Z(n402) );
  MUX21L U452 ( .A(n626), .B(n497), .S(n526), .Z(n401) );
  MUX21L U453 ( .A(n625), .B(n498), .S(n526), .Z(n400) );
  MUX21L U454 ( .A(n624), .B(n499), .S(n526), .Z(n399) );
  MUX21L U455 ( .A(n623), .B(n500), .S(n526), .Z(n398) );
  MUX21L U456 ( .A(n622), .B(n501), .S(n526), .Z(n397) );
  MUX21L U457 ( .A(n621), .B(n502), .S(n526), .Z(n396) );
  MUX21L U458 ( .A(n620), .B(n503), .S(n526), .Z(n395) );
  MUX21L U459 ( .A(n619), .B(n504), .S(n526), .Z(n394) );
  MUX21L U460 ( .A(n618), .B(n505), .S(n526), .Z(n393) );
  MUX21L U461 ( .A(n617), .B(n506), .S(n526), .Z(n392) );
  MUX21L U462 ( .A(n616), .B(n507), .S(n526), .Z(n391) );
  MUX21L U463 ( .A(n615), .B(n508), .S(n526), .Z(n390) );
  MUX21L U464 ( .A(n614), .B(n509), .S(n526), .Z(n389) );
  MUX21L U465 ( .A(n613), .B(n510), .S(n526), .Z(n388) );
  MUX21L U466 ( .A(n612), .B(n511), .S(n526), .Z(n387) );
  MUX21L U467 ( .A(n611), .B(n512), .S(n526), .Z(n386) );
  MUX21L U468 ( .A(n610), .B(n513), .S(n526), .Z(n385) );
  MUX21L U469 ( .A(n609), .B(n514), .S(n526), .Z(n384) );
  MUX21L U470 ( .A(n608), .B(n515), .S(n526), .Z(n383) );
  MUX21L U471 ( .A(n607), .B(n516), .S(n526), .Z(n382) );
  MUX21L U472 ( .A(n606), .B(n517), .S(n526), .Z(n381) );
  MUX21L U473 ( .A(n605), .B(n518), .S(n526), .Z(n380) );
  MUX21L U474 ( .A(n604), .B(n519), .S(n526), .Z(n379) );
  MUX21L U475 ( .A(n603), .B(n520), .S(n526), .Z(n378) );
  MUX21L U476 ( .A(n602), .B(n521), .S(n526), .Z(n377) );
  MUX21L U477 ( .A(n601), .B(n522), .S(n526), .Z(n376) );
  MUX21L U478 ( .A(n600), .B(n523), .S(n526), .Z(n375) );
  NR3 U479 ( .A(n524), .B(wr_ptr[0]), .C(n1), .Z(n526) );
  MUX21L U480 ( .A(n599), .B(n330), .S(n527), .Z(n374) );
  IV U481 ( .A(wr_data[0]), .Z(n330) );
  MUX21L U482 ( .A(n598), .B(n332), .S(n527), .Z(n373) );
  IV U483 ( .A(wr_data[35]), .Z(n332) );
  MUX21L U484 ( .A(n597), .B(n490), .S(n527), .Z(n372) );
  IV U485 ( .A(wr_data[34]), .Z(n490) );
  MUX21L U486 ( .A(n596), .B(n491), .S(n527), .Z(n371) );
  IV U487 ( .A(wr_data[33]), .Z(n491) );
  MUX21L U488 ( .A(n595), .B(n492), .S(n527), .Z(n370) );
  IV U489 ( .A(wr_data[32]), .Z(n492) );
  MUX21L U490 ( .A(n594), .B(n493), .S(n527), .Z(n369) );
  IV U491 ( .A(wr_data[31]), .Z(n493) );
  MUX21L U492 ( .A(n593), .B(n494), .S(n527), .Z(n368) );
  IV U493 ( .A(wr_data[30]), .Z(n494) );
  MUX21L U494 ( .A(n592), .B(n495), .S(n527), .Z(n367) );
  IV U495 ( .A(wr_data[29]), .Z(n495) );
  MUX21L U496 ( .A(n591), .B(n496), .S(n527), .Z(n366) );
  IV U497 ( .A(wr_data[28]), .Z(n496) );
  MUX21L U498 ( .A(n590), .B(n497), .S(n527), .Z(n365) );
  IV U499 ( .A(wr_data[27]), .Z(n497) );
  MUX21L U500 ( .A(n589), .B(n498), .S(n527), .Z(n364) );
  IV U501 ( .A(wr_data[26]), .Z(n498) );
  MUX21L U502 ( .A(n588), .B(n499), .S(n527), .Z(n363) );
  IV U503 ( .A(wr_data[25]), .Z(n499) );
  MUX21L U504 ( .A(n587), .B(n500), .S(n527), .Z(n362) );
  IV U505 ( .A(wr_data[24]), .Z(n500) );
  MUX21L U506 ( .A(n586), .B(n501), .S(n527), .Z(n361) );
  IV U507 ( .A(wr_data[23]), .Z(n501) );
  MUX21L U508 ( .A(n585), .B(n502), .S(n527), .Z(n360) );
  IV U509 ( .A(wr_data[22]), .Z(n502) );
  MUX21L U510 ( .A(n584), .B(n503), .S(n527), .Z(n359) );
  IV U511 ( .A(wr_data[21]), .Z(n503) );
  MUX21L U512 ( .A(n583), .B(n504), .S(n527), .Z(n358) );
  IV U513 ( .A(wr_data[20]), .Z(n504) );
  MUX21L U514 ( .A(n582), .B(n505), .S(n527), .Z(n357) );
  IV U515 ( .A(wr_data[19]), .Z(n505) );
  MUX21L U516 ( .A(n581), .B(n506), .S(n527), .Z(n356) );
  IV U517 ( .A(wr_data[18]), .Z(n506) );
  MUX21L U518 ( .A(n580), .B(n507), .S(n527), .Z(n355) );
  IV U519 ( .A(wr_data[17]), .Z(n507) );
  MUX21L U520 ( .A(n579), .B(n508), .S(n527), .Z(n354) );
  IV U521 ( .A(wr_data[16]), .Z(n508) );
  MUX21L U522 ( .A(n578), .B(n509), .S(n527), .Z(n353) );
  IV U523 ( .A(wr_data[15]), .Z(n509) );
  MUX21L U524 ( .A(n577), .B(n510), .S(n527), .Z(n352) );
  IV U525 ( .A(wr_data[14]), .Z(n510) );
  MUX21L U526 ( .A(n576), .B(n511), .S(n527), .Z(n351) );
  IV U527 ( .A(wr_data[13]), .Z(n511) );
  MUX21L U528 ( .A(n575), .B(n512), .S(n527), .Z(n350) );
  IV U529 ( .A(wr_data[12]), .Z(n512) );
  MUX21L U530 ( .A(n574), .B(n513), .S(n527), .Z(n349) );
  IV U531 ( .A(wr_data[11]), .Z(n513) );
  MUX21L U532 ( .A(n573), .B(n514), .S(n527), .Z(n348) );
  IV U533 ( .A(wr_data[10]), .Z(n514) );
  MUX21L U534 ( .A(n572), .B(n515), .S(n527), .Z(n347) );
  IV U535 ( .A(wr_data[9]), .Z(n515) );
  MUX21L U536 ( .A(n571), .B(n516), .S(n527), .Z(n346) );
  IV U537 ( .A(wr_data[8]), .Z(n516) );
  MUX21L U538 ( .A(n570), .B(n517), .S(n527), .Z(n345) );
  IV U539 ( .A(wr_data[7]), .Z(n517) );
  MUX21L U540 ( .A(n569), .B(n518), .S(n527), .Z(n344) );
  IV U541 ( .A(wr_data[6]), .Z(n518) );
  MUX21L U542 ( .A(n568), .B(n519), .S(n527), .Z(n343) );
  IV U543 ( .A(wr_data[5]), .Z(n519) );
  MUX21L U544 ( .A(n567), .B(n520), .S(n527), .Z(n342) );
  IV U545 ( .A(wr_data[4]), .Z(n520) );
  MUX21L U546 ( .A(n566), .B(n521), .S(n527), .Z(n341) );
  IV U547 ( .A(wr_data[3]), .Z(n521) );
  MUX21L U548 ( .A(n565), .B(n522), .S(n527), .Z(n340) );
  IV U549 ( .A(wr_data[2]), .Z(n522) );
  MUX21L U550 ( .A(n564), .B(n523), .S(n527), .Z(n339) );
  NR2 U551 ( .A(n528), .B(n524), .Z(n527) );
  IV U552 ( .A(wr_data[1]), .Z(n523) );
  AO7 U553 ( .A(wr_en), .B(n2), .C(n529), .Z(n338) );
  AO7 U554 ( .A(wr_en), .B(n563), .C(n529), .Z(n337) );
  AO7 U555 ( .A(n4), .B(n329), .C(n530), .Z(n336) );
  MUX21L U556 ( .A(grey_wr_ptr[0]), .B(n531), .S(wr_en), .Z(n530) );
  NR2 U557 ( .A(wr_ptr[0]), .B(n532), .Z(n531) );
  AO7 U558 ( .A(test_so4), .B(n329), .C(n533), .Z(n335) );
  EO1 U559 ( .A(grey_wr_ptr[1]), .B(n524), .C(n529), .D(n532), .Z(n533) );
  ND2 U560 ( .A(wr_en), .B(n534), .Z(n529) );
  EN U561 ( .A(test_so4), .B(n528), .Z(n534) );
  ND2 U562 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .Z(n528) );
  ND2 U563 ( .A(wr_en), .B(n532), .Z(n329) );
  EN U564 ( .A(n1), .B(wr_ptr[0]), .Z(n532) );
  AO4 U565 ( .A(n535), .B(n524), .C(n562), .D(n536), .Z(n334) );
  IV U566 ( .A(wr_en), .Z(n524) );
  AN2 U567 ( .A(n537), .B(n562), .Z(n535) );
  MUX21L U568 ( .A(n538), .B(n561), .S(n539), .Z(n333) );
  NR2 U569 ( .A(aempty), .B(n540), .Z(n539) );
  AO6 U570 ( .A(n541), .B(n542), .C(n561), .Z(n540) );
  IV U571 ( .A(rd_en), .Z(n538) );
  IV U572 ( .A(n537), .Z(afull) );
  AO3 U573 ( .A(n543), .B(n544), .C(n545), .D(n536), .Z(n537) );
  EO U574 ( .A(n546), .B(n547), .Z(n536) );
  EN U575 ( .A(sync_rd_ptr_1[2]), .B(n2), .Z(n547) );
  AO5 U576 ( .A(n544), .B(n548), .C(n1), .Z(n546) );
  EO U577 ( .A(sync_rd_ptr_1[2]), .B(sync_rd_ptr_1[1]), .Z(n548) );
  EO U578 ( .A(n549), .B(n550), .Z(n545) );
  EO U579 ( .A(wr_ptr[1]), .B(n544), .Z(n550) );
  NR2 U580 ( .A(wr_ptr[0]), .B(n551), .Z(n544) );
  AN2 U581 ( .A(wr_ptr[0]), .B(n551), .Z(n543) );
  EN U582 ( .A(n549), .B(sync_rd_ptr_1[0]), .Z(n551) );
  EN U583 ( .A(n711), .B(sync_rd_ptr_1[2]), .Z(n549) );
  IV U584 ( .A(n552), .Z(aempty) );
  AO3 U585 ( .A(n553), .B(n554), .C(n542), .D(n541), .Z(n552) );
  EO U586 ( .A(n555), .B(n556), .Z(n541) );
  NR2 U587 ( .A(n246), .B(n557), .Z(n556) );
  EN U588 ( .A(n712), .B(test_so5), .Z(n555) );
  EN U589 ( .A(n558), .B(n559), .Z(n542) );
  EO U590 ( .A(n557), .B(n246), .Z(n558) );
  IV U591 ( .A(n557), .Z(n554) );
  ND2 U592 ( .A(n560), .B(N45), .Z(n557) );
  NR2 U593 ( .A(n560), .B(N45), .Z(n553) );
  EN U594 ( .A(n559), .B(sync_wr_ptr_1_0_), .Z(n560) );
  EN U595 ( .A(n713), .B(test_so5), .Z(n559) );
endmodule

